// This is the unpowered netlist.
module cordic_tt_top (i_clk,
    i_rst_n,
    i_valid_in,
    o_valid_out,
    in_alpha,
    in_x,
    in_y,
    out_alpha,
    out_costheta,
    out_sintheta);
 input i_clk;
 input i_rst_n;
 input i_valid_in;
 output o_valid_out;
 input [17:0] in_alpha;
 input [17:0] in_x;
 input [17:0] in_y;
 output [17:0] out_alpha;
 output [17:0] out_costheta;
 output [17:0] out_sintheta;

 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.i_quadrant[0] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.i_quadrant[1] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[0] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[16] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[1] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ;
 wire \CORDIC_PE[0].genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[0] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[1] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[2] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[3] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[4] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[5] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[6] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[7] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[8] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[9] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[0] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[1] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[2] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[3] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[4] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[5] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[6] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[7] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ;
 wire \CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire clknet_0_i_clk;
 wire clknet_4_0_0_i_clk;
 wire clknet_4_10_0_i_clk;
 wire clknet_4_11_0_i_clk;
 wire clknet_4_12_0_i_clk;
 wire clknet_4_13_0_i_clk;
 wire clknet_4_14_0_i_clk;
 wire clknet_4_15_0_i_clk;
 wire clknet_4_1_0_i_clk;
 wire clknet_4_2_0_i_clk;
 wire clknet_4_3_0_i_clk;
 wire clknet_4_4_0_i_clk;
 wire clknet_4_5_0_i_clk;
 wire clknet_4_6_0_i_clk;
 wire clknet_4_7_0_i_clk;
 wire clknet_4_8_0_i_clk;
 wire clknet_4_9_0_i_clk;
 wire clknet_leaf_0_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_103_i_clk;
 wire clknet_leaf_104_i_clk;
 wire clknet_leaf_105_i_clk;
 wire clknet_leaf_106_i_clk;
 wire clknet_leaf_107_i_clk;
 wire clknet_leaf_108_i_clk;
 wire clknet_leaf_109_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_110_i_clk;
 wire clknet_leaf_111_i_clk;
 wire clknet_leaf_112_i_clk;
 wire clknet_leaf_113_i_clk;
 wire clknet_leaf_114_i_clk;
 wire clknet_leaf_115_i_clk;
 wire clknet_leaf_116_i_clk;
 wire clknet_leaf_117_i_clk;
 wire clknet_leaf_118_i_clk;
 wire clknet_leaf_119_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_120_i_clk;
 wire clknet_leaf_121_i_clk;
 wire clknet_leaf_122_i_clk;
 wire clknet_leaf_123_i_clk;
 wire clknet_leaf_124_i_clk;
 wire clknet_leaf_125_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_9_i_clk;
 wire \diff1[0] ;
 wire \diff1[10] ;
 wire \diff1[11] ;
 wire \diff1[12] ;
 wire \diff1[13] ;
 wire \diff1[14] ;
 wire \diff1[15] ;
 wire \diff1[16] ;
 wire \diff1[17] ;
 wire \diff1[1] ;
 wire \diff1[2] ;
 wire \diff1[3] ;
 wire \diff1[4] ;
 wire \diff1[5] ;
 wire \diff1[6] ;
 wire \diff1[7] ;
 wire \diff1[8] ;
 wire \diff1[9] ;
 wire \diff2[10] ;
 wire \diff2[11] ;
 wire \diff2[12] ;
 wire \diff2[13] ;
 wire \diff2[14] ;
 wire \diff2[15] ;
 wire \diff2[16] ;
 wire \diff2[17] ;
 wire \diff2[3] ;
 wire \diff2[4] ;
 wire \diff2[5] ;
 wire \diff2[6] ;
 wire \diff2[7] ;
 wire \diff2[8] ;
 wire \diff2[9] ;
 wire \diff3[10] ;
 wire \diff3[11] ;
 wire \diff3[12] ;
 wire \diff3[13] ;
 wire \diff3[14] ;
 wire \diff3[15] ;
 wire \diff3[16] ;
 wire \diff3[17] ;
 wire \diff3[4] ;
 wire \diff3[5] ;
 wire \diff3[6] ;
 wire \diff3[7] ;
 wire \diff3[8] ;
 wire \diff3[9] ;
 wire diff_valid;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \r_i_alpha1[10] ;
 wire \r_i_alpha1[11] ;
 wire \r_i_alpha1[12] ;
 wire \r_i_alpha1[13] ;
 wire \r_i_alpha1[14] ;
 wire \r_i_alpha1[15] ;
 wire \r_i_alpha1[16] ;
 wire \r_i_alpha1[17] ;
 wire \r_i_alpha1[4] ;
 wire \r_i_alpha1[5] ;
 wire \r_i_alpha1[6] ;
 wire \r_i_alpha1[7] ;
 wire \r_i_alpha1[8] ;
 wire \r_i_alpha1[9] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__buf_2 _07227_ (.A(net15),
    .X(_00991_));
 sky130_fd_sc_hd__clkbuf_4 _07228_ (.A(net2),
    .X(_00992_));
 sky130_fd_sc_hd__clkbuf_4 _07229_ (.A(_00992_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _07230_ (.A0(net365),
    .A1(_00991_),
    .S(_00993_),
    .X(_00994_));
 sky130_fd_sc_hd__clkbuf_1 _07231_ (.A(_00994_),
    .X(_00000_));
 sky130_fd_sc_hd__mux2_1 _07232_ (.A0(net332),
    .A1(net16),
    .S(_00993_),
    .X(_00995_));
 sky130_fd_sc_hd__clkbuf_1 _07233_ (.A(_00995_),
    .X(_00001_));
 sky130_fd_sc_hd__mux2_1 _07234_ (.A0(net353),
    .A1(net17),
    .S(_00993_),
    .X(_00996_));
 sky130_fd_sc_hd__clkbuf_1 _07235_ (.A(_00996_),
    .X(_00002_));
 sky130_fd_sc_hd__mux2_1 _07236_ (.A0(net341),
    .A1(net18),
    .S(_00993_),
    .X(_00997_));
 sky130_fd_sc_hd__clkbuf_1 _07237_ (.A(_00997_),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _07238_ (.A0(net368),
    .A1(net19),
    .S(_00993_),
    .X(_00998_));
 sky130_fd_sc_hd__clkbuf_1 _07239_ (.A(_00998_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _07240_ (.A0(net329),
    .A1(net20),
    .S(_00993_),
    .X(_00999_));
 sky130_fd_sc_hd__clkbuf_1 _07241_ (.A(_00999_),
    .X(_00005_));
 sky130_fd_sc_hd__buf_4 _07242_ (.A(_00992_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _07243_ (.A0(net344),
    .A1(net4),
    .S(_01000_),
    .X(_01001_));
 sky130_fd_sc_hd__clkbuf_1 _07244_ (.A(_01001_),
    .X(_00006_));
 sky130_fd_sc_hd__mux2_1 _07245_ (.A0(net338),
    .A1(net5),
    .S(_01000_),
    .X(_01002_));
 sky130_fd_sc_hd__clkbuf_1 _07246_ (.A(_01002_),
    .X(_00007_));
 sky130_fd_sc_hd__clkbuf_4 _07247_ (.A(net6),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _07248_ (.A0(net367),
    .A1(_01003_),
    .S(_01000_),
    .X(_01004_));
 sky130_fd_sc_hd__clkbuf_1 _07249_ (.A(_01004_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _07250_ (.A0(net354),
    .A1(net7),
    .S(_01000_),
    .X(_01005_));
 sky130_fd_sc_hd__clkbuf_1 _07251_ (.A(_01005_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _07252_ (.A0(net363),
    .A1(net8),
    .S(_01000_),
    .X(_01006_));
 sky130_fd_sc_hd__clkbuf_1 _07253_ (.A(_01006_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _07254_ (.A0(net386),
    .A1(net9),
    .S(_01000_),
    .X(_01007_));
 sky130_fd_sc_hd__clkbuf_1 _07255_ (.A(_01007_),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _07256_ (.A0(net376),
    .A1(net10),
    .S(_01000_),
    .X(_01008_));
 sky130_fd_sc_hd__clkbuf_1 _07257_ (.A(_01008_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _07258_ (.A0(net178),
    .A1(net11),
    .S(_01000_),
    .X(_01009_));
 sky130_fd_sc_hd__clkbuf_1 _07259_ (.A(_01009_),
    .X(_00013_));
 sky130_fd_sc_hd__buf_2 _07260_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _07261_ (.A0(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .S(_01010_),
    .X(_01011_));
 sky130_fd_sc_hd__buf_4 _07262_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_01012_));
 sky130_fd_sc_hd__buf_4 _07263_ (.A(_01012_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _07264_ (.A0(net385),
    .A1(_01011_),
    .S(_01013_),
    .X(_01014_));
 sky130_fd_sc_hd__clkbuf_1 _07265_ (.A(_01014_),
    .X(_00014_));
 sky130_fd_sc_hd__inv_2 _07266_ (.A(_01012_),
    .Y(_01015_));
 sky130_fd_sc_hd__clkbuf_4 _07267_ (.A(_01015_),
    .X(_01016_));
 sky130_fd_sc_hd__inv_2 _07268_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .Y(_01017_));
 sky130_fd_sc_hd__or2_1 _07269_ (.A(_01017_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(_01018_));
 sky130_fd_sc_hd__buf_2 _07270_ (.A(_01018_),
    .X(_01019_));
 sky130_fd_sc_hd__xnor2_1 _07271_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_01020_));
 sky130_fd_sc_hd__inv_2 _07272_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .Y(_01021_));
 sky130_fd_sc_hd__clkbuf_4 _07273_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(_01022_));
 sky130_fd_sc_hd__nand2_1 _07274_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_01010_),
    .Y(_01023_));
 sky130_fd_sc_hd__xnor2_1 _07275_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .Y(_01024_));
 sky130_fd_sc_hd__or2_1 _07276_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(_01025_));
 sky130_fd_sc_hd__buf_2 _07277_ (.A(_01025_),
    .X(_01026_));
 sky130_fd_sc_hd__o221a_1 _07278_ (.A1(_01021_),
    .A2(_01022_),
    .B1(_01023_),
    .B2(_01024_),
    .C1(_01026_),
    .X(_01027_));
 sky130_fd_sc_hd__o21ai_1 _07279_ (.A1(_01019_),
    .A2(_01020_),
    .B1(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__clkbuf_4 _07280_ (.A(_01026_),
    .X(_01029_));
 sky130_fd_sc_hd__clkbuf_4 _07281_ (.A(_01012_),
    .X(_01030_));
 sky130_fd_sc_hd__o21a_1 _07282_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .A2(_01029_),
    .B1(_01030_),
    .X(_01031_));
 sky130_fd_sc_hd__a22o_1 _07283_ (.A1(_01016_),
    .A2(net243),
    .B1(_01028_),
    .B2(_01031_),
    .X(_00015_));
 sky130_fd_sc_hd__inv_2 _07284_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_01032_));
 sky130_fd_sc_hd__or3_1 _07285_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .C(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(_01033_));
 sky130_fd_sc_hd__o21ai_1 _07286_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _07287_ (.A(_01033_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__o221a_1 _07288_ (.A1(_01032_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B1(_01019_),
    .B2(_01035_),
    .C1(_01026_),
    .X(_01036_));
 sky130_fd_sc_hd__and2_1 _07289_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_01010_),
    .X(_01037_));
 sky130_fd_sc_hd__or3_4 _07290_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .C(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(_01038_));
 sky130_fd_sc_hd__o21ai_1 _07291_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_01039_));
 sky130_fd_sc_hd__and2_1 _07292_ (.A(_01038_),
    .B(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__nand2_1 _07293_ (.A(_01037_),
    .B(_01040_),
    .Y(_01041_));
 sky130_fd_sc_hd__o2bb2a_1 _07294_ (.A1_N(_01036_),
    .A2_N(_01041_),
    .B1(_01026_),
    .B2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _07295_ (.A0(net370),
    .A1(_01042_),
    .S(_01013_),
    .X(_01043_));
 sky130_fd_sc_hd__clkbuf_1 _07296_ (.A(_01043_),
    .X(_00016_));
 sky130_fd_sc_hd__clkbuf_4 _07297_ (.A(_01015_),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_4 _07298_ (.A(_01026_),
    .X(_01045_));
 sky130_fd_sc_hd__nor2_1 _07299_ (.A(_01017_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .Y(_01046_));
 sky130_fd_sc_hd__buf_2 _07300_ (.A(_01046_),
    .X(_01047_));
 sky130_fd_sc_hd__or4_4 _07301_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .C(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .D(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(_01048_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_01033_),
    .Y(_01049_));
 sky130_fd_sc_hd__and3_1 _07303_ (.A(_01047_),
    .B(_01048_),
    .C(_01049_),
    .X(_01050_));
 sky130_fd_sc_hd__clkbuf_4 _07304_ (.A(_01017_),
    .X(_01051_));
 sky130_fd_sc_hd__clkbuf_4 _07305_ (.A(_01037_),
    .X(_01052_));
 sky130_fd_sc_hd__or2_1 _07306_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_01038_),
    .X(_01053_));
 sky130_fd_sc_hd__nand2_1 _07307_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_01038_),
    .Y(_01054_));
 sky130_fd_sc_hd__and2_1 _07308_ (.A(_01053_),
    .B(_01054_),
    .X(_01055_));
 sky130_fd_sc_hd__nor2_1 _07309_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_01010_),
    .Y(_01056_));
 sky130_fd_sc_hd__clkbuf_4 _07310_ (.A(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__a221o_1 _07311_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01055_),
    .C1(_01057_),
    .X(_01058_));
 sky130_fd_sc_hd__buf_4 _07312_ (.A(_01012_),
    .X(_01059_));
 sky130_fd_sc_hd__o221a_1 _07313_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A2(_01045_),
    .B1(_01050_),
    .B2(_01058_),
    .C1(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__a21o_1 _07314_ (.A1(_01044_),
    .A2(net171),
    .B1(_01060_),
    .X(_00017_));
 sky130_fd_sc_hd__xnor2_1 _07315_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_01048_),
    .Y(_01061_));
 sky130_fd_sc_hd__nor2_1 _07316_ (.A(_01019_),
    .B(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__xor2_1 _07317_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_01053_),
    .X(_01063_));
 sky130_fd_sc_hd__a221o_1 _07318_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01063_),
    .C1(_01057_),
    .X(_01064_));
 sky130_fd_sc_hd__o221a_1 _07319_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(_01045_),
    .B1(_01062_),
    .B2(_01064_),
    .C1(_01059_),
    .X(_01065_));
 sky130_fd_sc_hd__a21o_1 _07320_ (.A1(_01044_),
    .A2(net168),
    .B1(_01065_),
    .X(_00018_));
 sky130_fd_sc_hd__or3_4 _07321_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .C(_01048_),
    .X(_01066_));
 sky130_fd_sc_hd__o21ai_1 _07322_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(_01048_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .Y(_01067_));
 sky130_fd_sc_hd__and3_1 _07323_ (.A(_01047_),
    .B(_01066_),
    .C(_01067_),
    .X(_01068_));
 sky130_fd_sc_hd__or4_4 _07324_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .C(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .D(_01038_),
    .X(_01069_));
 sky130_fd_sc_hd__o21ai_1 _07325_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A2(_01053_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .Y(_01070_));
 sky130_fd_sc_hd__and2_1 _07326_ (.A(_01069_),
    .B(_01070_),
    .X(_01071_));
 sky130_fd_sc_hd__clkbuf_4 _07327_ (.A(_01056_),
    .X(_01072_));
 sky130_fd_sc_hd__a221o_1 _07328_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(_01017_),
    .B1(_01052_),
    .B2(_01071_),
    .C1(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__or2_1 _07329_ (.A(_01068_),
    .B(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__o21a_1 _07330_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_01029_),
    .B1(_01030_),
    .X(_01075_));
 sky130_fd_sc_hd__a22o_1 _07331_ (.A1(_01016_),
    .A2(net284),
    .B1(_01074_),
    .B2(_01075_),
    .X(_00019_));
 sky130_fd_sc_hd__clkbuf_4 _07332_ (.A(_01046_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_4 _07333_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_01066_),
    .X(_01077_));
 sky130_fd_sc_hd__nand2_1 _07334_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_01066_),
    .Y(_01078_));
 sky130_fd_sc_hd__and2_1 _07335_ (.A(_01077_),
    .B(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__buf_2 _07336_ (.A(_01017_),
    .X(_01080_));
 sky130_fd_sc_hd__clkbuf_4 _07337_ (.A(_01037_),
    .X(_01081_));
 sky130_fd_sc_hd__or2_4 _07338_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_01069_),
    .X(_01082_));
 sky130_fd_sc_hd__nand2_1 _07339_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_01069_),
    .Y(_01083_));
 sky130_fd_sc_hd__and2_1 _07340_ (.A(_01082_),
    .B(_01083_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_4 _07341_ (.A(_01056_),
    .X(_01085_));
 sky130_fd_sc_hd__a221o_1 _07342_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A2(_01080_),
    .B1(_01081_),
    .B2(_01084_),
    .C1(_01085_),
    .X(_01086_));
 sky130_fd_sc_hd__a21o_1 _07343_ (.A1(_01076_),
    .A2(_01079_),
    .B1(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__clkbuf_4 _07344_ (.A(_01012_),
    .X(_01088_));
 sky130_fd_sc_hd__o21a_1 _07345_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01089_));
 sky130_fd_sc_hd__a22o_1 _07346_ (.A1(_01016_),
    .A2(net279),
    .B1(_01087_),
    .B2(_01089_),
    .X(_00020_));
 sky130_fd_sc_hd__xnor2_1 _07347_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_01077_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _07348_ (.A(_01019_),
    .B(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__xor2_1 _07349_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_01082_),
    .X(_01092_));
 sky130_fd_sc_hd__a221o_1 _07350_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01092_),
    .C1(_01057_),
    .X(_01093_));
 sky130_fd_sc_hd__o221a_1 _07351_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(_01045_),
    .B1(_01091_),
    .B2(_01093_),
    .C1(_01059_),
    .X(_01094_));
 sky130_fd_sc_hd__a21o_1 _07352_ (.A1(_01044_),
    .A2(net185),
    .B1(_01094_),
    .X(_00021_));
 sky130_fd_sc_hd__clkbuf_4 _07353_ (.A(_01015_),
    .X(_01095_));
 sky130_fd_sc_hd__or3_1 _07354_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .C(_01077_),
    .X(_01096_));
 sky130_fd_sc_hd__o21ai_1 _07355_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(_01077_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .Y(_01097_));
 sky130_fd_sc_hd__and3_1 _07356_ (.A(_01047_),
    .B(_01096_),
    .C(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__or3_1 _07357_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .C(_01082_),
    .X(_01099_));
 sky130_fd_sc_hd__o21ai_1 _07358_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(_01082_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_01100_));
 sky130_fd_sc_hd__and2_1 _07359_ (.A(_01099_),
    .B(_01100_),
    .X(_01101_));
 sky130_fd_sc_hd__a221o_1 _07360_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_01017_),
    .B1(_01052_),
    .B2(_01101_),
    .C1(_01072_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _07361_ (.A(_01098_),
    .B(_01102_),
    .X(_01103_));
 sky130_fd_sc_hd__o21a_1 _07362_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01104_));
 sky130_fd_sc_hd__a22o_1 _07363_ (.A1(_01095_),
    .A2(net233),
    .B1(_01103_),
    .B2(_01104_),
    .X(_00022_));
 sky130_fd_sc_hd__or2_4 _07364_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_01096_),
    .X(_01105_));
 sky130_fd_sc_hd__nand2_1 _07365_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_01096_),
    .Y(_01106_));
 sky130_fd_sc_hd__and2_1 _07366_ (.A(_01105_),
    .B(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_4 _07367_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_01099_),
    .X(_01108_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_01099_),
    .Y(_01109_));
 sky130_fd_sc_hd__and2_1 _07369_ (.A(_01108_),
    .B(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__a221o_1 _07370_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_01080_),
    .B1(_01081_),
    .B2(_01110_),
    .C1(_01085_),
    .X(_01111_));
 sky130_fd_sc_hd__a21o_1 _07371_ (.A1(_01076_),
    .A2(_01107_),
    .B1(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__o21a_1 _07372_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01113_));
 sky130_fd_sc_hd__a22o_1 _07373_ (.A1(_01095_),
    .A2(net208),
    .B1(_01112_),
    .B2(_01113_),
    .X(_00023_));
 sky130_fd_sc_hd__xnor2_1 _07374_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_01105_),
    .Y(_01114_));
 sky130_fd_sc_hd__nor2_1 _07375_ (.A(_01019_),
    .B(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__xor2_1 _07376_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_01108_),
    .X(_01116_));
 sky130_fd_sc_hd__a221o_1 _07377_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01116_),
    .C1(_01057_),
    .X(_01117_));
 sky130_fd_sc_hd__o221a_1 _07378_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_01045_),
    .B1(_01115_),
    .B2(_01117_),
    .C1(_01059_),
    .X(_01118_));
 sky130_fd_sc_hd__a21o_1 _07379_ (.A1(_01044_),
    .A2(net182),
    .B1(_01118_),
    .X(_00024_));
 sky130_fd_sc_hd__or3_4 _07380_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .C(_01105_),
    .X(_01119_));
 sky130_fd_sc_hd__o21ai_1 _07381_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_01105_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .Y(_01120_));
 sky130_fd_sc_hd__and3_1 _07382_ (.A(_01047_),
    .B(_01119_),
    .C(_01120_),
    .X(_01121_));
 sky130_fd_sc_hd__clkbuf_4 _07383_ (.A(_01037_),
    .X(_01122_));
 sky130_fd_sc_hd__or3_1 _07384_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .C(_01108_),
    .X(_01123_));
 sky130_fd_sc_hd__o21ai_1 _07385_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_01108_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .Y(_01124_));
 sky130_fd_sc_hd__and2_1 _07386_ (.A(_01123_),
    .B(_01124_),
    .X(_01125_));
 sky130_fd_sc_hd__a221o_1 _07387_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_01017_),
    .B1(_01122_),
    .B2(_01125_),
    .C1(_01072_),
    .X(_01126_));
 sky130_fd_sc_hd__or2_1 _07388_ (.A(_01121_),
    .B(_01126_),
    .X(_01127_));
 sky130_fd_sc_hd__o21a_1 _07389_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01128_));
 sky130_fd_sc_hd__a22o_1 _07390_ (.A1(_01095_),
    .A2(net230),
    .B1(_01127_),
    .B2(_01128_),
    .X(_00025_));
 sky130_fd_sc_hd__or2_1 _07391_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_01119_),
    .X(_01129_));
 sky130_fd_sc_hd__nand2_1 _07392_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_01119_),
    .Y(_01130_));
 sky130_fd_sc_hd__and2_1 _07393_ (.A(_01129_),
    .B(_01130_),
    .X(_01131_));
 sky130_fd_sc_hd__or2_4 _07394_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_01123_),
    .X(_01132_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_01123_),
    .Y(_01133_));
 sky130_fd_sc_hd__and2_1 _07396_ (.A(_01132_),
    .B(_01133_),
    .X(_01134_));
 sky130_fd_sc_hd__a221o_1 _07397_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_01080_),
    .B1(_01081_),
    .B2(_01134_),
    .C1(_01085_),
    .X(_01135_));
 sky130_fd_sc_hd__a21o_1 _07398_ (.A1(_01076_),
    .A2(_01131_),
    .B1(_01135_),
    .X(_01136_));
 sky130_fd_sc_hd__o21a_1 _07399_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01137_));
 sky130_fd_sc_hd__a22o_1 _07400_ (.A1(_01095_),
    .A2(net197),
    .B1(_01136_),
    .B2(_01137_),
    .X(_00026_));
 sky130_fd_sc_hd__xnor2_1 _07401_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_01129_),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_1 _07402_ (.A(_01019_),
    .B(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__xor2_1 _07403_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_01132_),
    .X(_01140_));
 sky130_fd_sc_hd__a221o_1 _07404_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01140_),
    .C1(_01057_),
    .X(_01141_));
 sky130_fd_sc_hd__o221a_1 _07405_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_01045_),
    .B1(_01139_),
    .B2(_01141_),
    .C1(_01059_),
    .X(_01142_));
 sky130_fd_sc_hd__a21o_1 _07406_ (.A1(_01044_),
    .A2(net170),
    .B1(_01142_),
    .X(_00027_));
 sky130_fd_sc_hd__or3_4 _07407_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .C(_01129_),
    .X(_01143_));
 sky130_fd_sc_hd__o21ai_1 _07408_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_01129_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .Y(_01144_));
 sky130_fd_sc_hd__and2_1 _07409_ (.A(_01143_),
    .B(_01144_),
    .X(_01145_));
 sky130_fd_sc_hd__or3_1 _07410_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .C(_01132_),
    .X(_01146_));
 sky130_fd_sc_hd__o21ai_1 _07411_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_01132_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .Y(_01147_));
 sky130_fd_sc_hd__and2_1 _07412_ (.A(_01146_),
    .B(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__a221o_1 _07413_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_01051_),
    .B1(_01081_),
    .B2(_01148_),
    .C1(_01085_),
    .X(_01149_));
 sky130_fd_sc_hd__a21o_1 _07414_ (.A1(_01076_),
    .A2(_01145_),
    .B1(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__o21a_1 _07415_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01151_));
 sky130_fd_sc_hd__a22o_1 _07416_ (.A1(_01095_),
    .A2(net249),
    .B1(_01150_),
    .B2(_01151_),
    .X(_00028_));
 sky130_fd_sc_hd__xnor2_1 _07417_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_01143_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _07418_ (.A(_01019_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__or2_1 _07419_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_01146_),
    .X(_01154_));
 sky130_fd_sc_hd__nand2_1 _07420_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_01146_),
    .Y(_01155_));
 sky130_fd_sc_hd__and2_1 _07421_ (.A(_01154_),
    .B(_01155_),
    .X(_01156_));
 sky130_fd_sc_hd__a221o_1 _07422_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01156_),
    .C1(_01057_),
    .X(_01157_));
 sky130_fd_sc_hd__o221a_1 _07423_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_01045_),
    .B1(_01153_),
    .B2(_01157_),
    .C1(_01059_),
    .X(_01158_));
 sky130_fd_sc_hd__a21o_1 _07424_ (.A1(_01044_),
    .A2(net177),
    .B1(_01158_),
    .X(_00029_));
 sky130_fd_sc_hd__clkbuf_4 _07425_ (.A(_01026_),
    .X(_01159_));
 sky130_fd_sc_hd__or2_1 _07426_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_01143_),
    .X(_01160_));
 sky130_fd_sc_hd__or2_1 _07427_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__nand2_1 _07428_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_01160_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _07429_ (.A(_01161_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _07430_ (.A(_01019_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__nor2_2 _07431_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_01154_),
    .Y(_01165_));
 sky130_fd_sc_hd__and2_1 _07432_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_01154_),
    .X(_01166_));
 sky130_fd_sc_hd__nor2_1 _07433_ (.A(_01165_),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__a221o_1 _07434_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_01051_),
    .B1(_01052_),
    .B2(_01167_),
    .C1(_01057_),
    .X(_01168_));
 sky130_fd_sc_hd__o221a_1 _07435_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(_01159_),
    .B1(_01164_),
    .B2(_01168_),
    .C1(_01059_),
    .X(_01169_));
 sky130_fd_sc_hd__a21o_1 _07436_ (.A1(_01044_),
    .A2(net193),
    .B1(_01169_),
    .X(_00030_));
 sky130_fd_sc_hd__xnor2_1 _07437_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_01161_),
    .Y(_01170_));
 sky130_fd_sc_hd__inv_2 _07438_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_01171_));
 sky130_fd_sc_hd__xnor2_1 _07439_ (.A(_01171_),
    .B(_01165_),
    .Y(_01172_));
 sky130_fd_sc_hd__o221a_1 _07440_ (.A1(_01171_),
    .A2(_01022_),
    .B1(_01023_),
    .B2(_01172_),
    .C1(_01026_),
    .X(_01173_));
 sky130_fd_sc_hd__o21ai_1 _07441_ (.A1(_01019_),
    .A2(_01170_),
    .B1(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__o21a_1 _07442_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01175_));
 sky130_fd_sc_hd__a22o_1 _07443_ (.A1(_01095_),
    .A2(net306),
    .B1(_01174_),
    .B2(_01175_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _07444_ (.A0(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .S(_01010_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _07445_ (.A0(net76),
    .A1(_01176_),
    .S(_01013_),
    .X(_01177_));
 sky130_fd_sc_hd__clkbuf_1 _07446_ (.A(_01177_),
    .X(_00032_));
 sky130_fd_sc_hd__a2bb2o_1 _07447_ (.A1_N(_01010_),
    .A2_N(_01024_),
    .B1(_01052_),
    .B2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_01178_));
 sky130_fd_sc_hd__a21oi_1 _07448_ (.A1(_01010_),
    .A2(_01020_),
    .B1(_01022_),
    .Y(_01179_));
 sky130_fd_sc_hd__o221a_1 _07449_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .A2(_01159_),
    .B1(_01178_),
    .B2(_01179_),
    .C1(_01059_),
    .X(_01180_));
 sky130_fd_sc_hd__a21o_1 _07450_ (.A1(_01044_),
    .A2(net439),
    .B1(_01180_),
    .X(_00033_));
 sky130_fd_sc_hd__a32o_1 _07451_ (.A1(_01051_),
    .A2(_01033_),
    .A3(_01034_),
    .B1(_01081_),
    .B2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .X(_01181_));
 sky130_fd_sc_hd__a211o_1 _07452_ (.A1(_01076_),
    .A2(_01040_),
    .B1(_01181_),
    .C1(_01085_),
    .X(_01182_));
 sky130_fd_sc_hd__a21oi_1 _07453_ (.A1(_01032_),
    .A2(_01085_),
    .B1(_01015_),
    .Y(_01183_));
 sky130_fd_sc_hd__a22o_1 _07454_ (.A1(_01095_),
    .A2(net617),
    .B1(_01182_),
    .B2(_01183_),
    .X(_00034_));
 sky130_fd_sc_hd__a32o_1 _07455_ (.A1(_01051_),
    .A2(_01048_),
    .A3(_01049_),
    .B1(_01076_),
    .B2(_01055_),
    .X(_01184_));
 sky130_fd_sc_hd__a211o_1 _07456_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A2(_01081_),
    .B1(_01184_),
    .C1(_01085_),
    .X(_01185_));
 sky130_fd_sc_hd__o21a_1 _07457_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A2(_01029_),
    .B1(_01088_),
    .X(_01186_));
 sky130_fd_sc_hd__a22o_1 _07458_ (.A1(_01095_),
    .A2(net609),
    .B1(_01185_),
    .B2(_01186_),
    .X(_00035_));
 sky130_fd_sc_hd__nor2_1 _07459_ (.A(_01022_),
    .B(_01061_),
    .Y(_01187_));
 sky130_fd_sc_hd__a221o_1 _07460_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(_01122_),
    .B1(_01063_),
    .B2(_01047_),
    .C1(_01057_),
    .X(_01188_));
 sky130_fd_sc_hd__o221a_1 _07461_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A2(_01159_),
    .B1(_01187_),
    .B2(_01188_),
    .C1(_01059_),
    .X(_01189_));
 sky130_fd_sc_hd__a21o_1 _07462_ (.A1(_01044_),
    .A2(net374),
    .B1(_01189_),
    .X(_00036_));
 sky130_fd_sc_hd__and3_1 _07463_ (.A(_01080_),
    .B(_01066_),
    .C(_01067_),
    .X(_01190_));
 sky130_fd_sc_hd__a221o_1 _07464_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_01122_),
    .B1(_01071_),
    .B2(_01047_),
    .C1(_01057_),
    .X(_01191_));
 sky130_fd_sc_hd__o221a_1 _07465_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(_01159_),
    .B1(_01190_),
    .B2(_01191_),
    .C1(_01030_),
    .X(_01192_));
 sky130_fd_sc_hd__a21o_1 _07466_ (.A1(_01044_),
    .A2(net335),
    .B1(_01192_),
    .X(_00037_));
 sky130_fd_sc_hd__a21o_1 _07467_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(_01081_),
    .B1(_01085_),
    .X(_01193_));
 sky130_fd_sc_hd__a221o_1 _07468_ (.A1(_01076_),
    .A2(_01084_),
    .B1(_01079_),
    .B2(_01080_),
    .C1(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__o21a_1 _07469_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A2(_01045_),
    .B1(_01088_),
    .X(_01195_));
 sky130_fd_sc_hd__a22o_1 _07470_ (.A1(_01095_),
    .A2(net452),
    .B1(_01194_),
    .B2(_01195_),
    .X(_00038_));
 sky130_fd_sc_hd__nor2_1 _07471_ (.A(_01022_),
    .B(_01090_),
    .Y(_01196_));
 sky130_fd_sc_hd__a221o_1 _07472_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(_01122_),
    .B1(_01092_),
    .B2(_01047_),
    .C1(_01072_),
    .X(_01197_));
 sky130_fd_sc_hd__o221a_1 _07473_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(_01159_),
    .B1(_01196_),
    .B2(_01197_),
    .C1(_01030_),
    .X(_01198_));
 sky130_fd_sc_hd__a21o_1 _07474_ (.A1(_01016_),
    .A2(net328),
    .B1(_01198_),
    .X(_00039_));
 sky130_fd_sc_hd__and3_1 _07475_ (.A(_01080_),
    .B(_01096_),
    .C(_01097_),
    .X(_01199_));
 sky130_fd_sc_hd__a221o_1 _07476_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_01122_),
    .B1(_01101_),
    .B2(_01047_),
    .C1(_01072_),
    .X(_01200_));
 sky130_fd_sc_hd__o221a_1 _07477_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_01159_),
    .B1(_01199_),
    .B2(_01200_),
    .C1(_01030_),
    .X(_01201_));
 sky130_fd_sc_hd__a21o_1 _07478_ (.A1(_01016_),
    .A2(net302),
    .B1(_01201_),
    .X(_00040_));
 sky130_fd_sc_hd__a21o_1 _07479_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_01081_),
    .B1(_01085_),
    .X(_01202_));
 sky130_fd_sc_hd__a221o_1 _07480_ (.A1(_01076_),
    .A2(_01110_),
    .B1(_01107_),
    .B2(_01080_),
    .C1(_01202_),
    .X(_01203_));
 sky130_fd_sc_hd__o21a_1 _07481_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_01045_),
    .B1(_01088_),
    .X(_01204_));
 sky130_fd_sc_hd__a22o_1 _07482_ (.A1(_01095_),
    .A2(net369),
    .B1(_01203_),
    .B2(_01204_),
    .X(_00041_));
 sky130_fd_sc_hd__nor2_1 _07483_ (.A(_01022_),
    .B(_01114_),
    .Y(_01205_));
 sky130_fd_sc_hd__a221o_1 _07484_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_01122_),
    .B1(_01116_),
    .B2(_01047_),
    .C1(_01072_),
    .X(_01206_));
 sky130_fd_sc_hd__o221a_1 _07485_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_01159_),
    .B1(_01205_),
    .B2(_01206_),
    .C1(_01030_),
    .X(_01207_));
 sky130_fd_sc_hd__a21o_1 _07486_ (.A1(_01016_),
    .A2(net253),
    .B1(_01207_),
    .X(_00042_));
 sky130_fd_sc_hd__and3_1 _07487_ (.A(_01080_),
    .B(_01119_),
    .C(_01120_),
    .X(_01208_));
 sky130_fd_sc_hd__a221o_1 _07488_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_01122_),
    .B1(_01125_),
    .B2(_01047_),
    .C1(_01072_),
    .X(_01209_));
 sky130_fd_sc_hd__o221a_1 _07489_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_01159_),
    .B1(_01208_),
    .B2(_01209_),
    .C1(_01030_),
    .X(_01210_));
 sky130_fd_sc_hd__a21o_1 _07490_ (.A1(_01016_),
    .A2(net255),
    .B1(_01210_),
    .X(_00043_));
 sky130_fd_sc_hd__a21o_1 _07491_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_01081_),
    .B1(_01085_),
    .X(_01211_));
 sky130_fd_sc_hd__a221o_1 _07492_ (.A1(_01076_),
    .A2(_01134_),
    .B1(_01131_),
    .B2(_01080_),
    .C1(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__o21a_1 _07493_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_01045_),
    .B1(_01013_),
    .X(_01213_));
 sky130_fd_sc_hd__a22o_1 _07494_ (.A1(_01015_),
    .A2(net505),
    .B1(_01212_),
    .B2(_01213_),
    .X(_00044_));
 sky130_fd_sc_hd__nor2_1 _07495_ (.A(_01022_),
    .B(_01138_),
    .Y(_01214_));
 sky130_fd_sc_hd__a221o_1 _07496_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_01122_),
    .B1(_01140_),
    .B2(_01046_),
    .C1(_01072_),
    .X(_01215_));
 sky130_fd_sc_hd__o221a_1 _07497_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_01159_),
    .B1(_01214_),
    .B2(_01215_),
    .C1(_01030_),
    .X(_01216_));
 sky130_fd_sc_hd__a21o_1 _07498_ (.A1(_01016_),
    .A2(net231),
    .B1(_01216_),
    .X(_00045_));
 sky130_fd_sc_hd__a21o_1 _07499_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_01081_),
    .B1(_01057_),
    .X(_01217_));
 sky130_fd_sc_hd__a221o_1 _07500_ (.A1(_01076_),
    .A2(_01148_),
    .B1(_01145_),
    .B2(_01080_),
    .C1(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__o21a_1 _07501_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_01045_),
    .B1(_01013_),
    .X(_01219_));
 sky130_fd_sc_hd__a22o_1 _07502_ (.A1(_01015_),
    .A2(net477),
    .B1(_01218_),
    .B2(_01219_),
    .X(_00046_));
 sky130_fd_sc_hd__nor2_1 _07503_ (.A(_01022_),
    .B(_01152_),
    .Y(_01220_));
 sky130_fd_sc_hd__a221o_1 _07504_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_01122_),
    .B1(_01156_),
    .B2(_01046_),
    .C1(_01072_),
    .X(_01221_));
 sky130_fd_sc_hd__o221a_1 _07505_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(_01159_),
    .B1(_01220_),
    .B2(_01221_),
    .C1(_01030_),
    .X(_01222_));
 sky130_fd_sc_hd__a21o_1 _07506_ (.A1(_01016_),
    .A2(net214),
    .B1(_01222_),
    .X(_00047_));
 sky130_fd_sc_hd__nor2_1 _07507_ (.A(_01022_),
    .B(_01163_),
    .Y(_01223_));
 sky130_fd_sc_hd__a221o_1 _07508_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(_01122_),
    .B1(_01167_),
    .B2(_01046_),
    .C1(_01072_),
    .X(_01224_));
 sky130_fd_sc_hd__o221a_1 _07509_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_01026_),
    .B1(_01223_),
    .B2(_01224_),
    .C1(_01030_),
    .X(_01225_));
 sky130_fd_sc_hd__a21o_1 _07510_ (.A1(_01016_),
    .A2(net229),
    .B1(_01225_),
    .X(_00048_));
 sky130_fd_sc_hd__a21oi_1 _07511_ (.A1(_01010_),
    .A2(_01170_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .Y(_01226_));
 sky130_fd_sc_hd__a2bb2o_1 _07512_ (.A1_N(_01010_),
    .A2_N(_01172_),
    .B1(_01037_),
    .B2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_01227_));
 sky130_fd_sc_hd__o22a_1 _07513_ (.A1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_01026_),
    .B1(_01226_),
    .B2(_01227_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _07514_ (.A0(net416),
    .A1(_01228_),
    .S(_01013_),
    .X(_01229_));
 sky130_fd_sc_hd__clkbuf_1 _07515_ (.A(_01229_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _07516_ (.A0(net371),
    .A1(net245),
    .S(_01013_),
    .X(_01230_));
 sky130_fd_sc_hd__clkbuf_1 _07517_ (.A(_01230_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _07518_ (.A0(net67),
    .A1(net318),
    .S(_01013_),
    .X(_01231_));
 sky130_fd_sc_hd__clkbuf_1 _07519_ (.A(net319),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _07520_ (.A0(net421),
    .A1(net323),
    .S(_01013_),
    .X(_01232_));
 sky130_fd_sc_hd__clkbuf_1 _07521_ (.A(_01232_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _07522_ (.A0(net69),
    .A1(net303),
    .S(_01013_),
    .X(_01233_));
 sky130_fd_sc_hd__clkbuf_1 _07523_ (.A(net304),
    .X(_00053_));
 sky130_fd_sc_hd__clkbuf_4 _07524_ (.A(_01012_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _07525_ (.A0(net373),
    .A1(net316),
    .S(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__clkbuf_1 _07526_ (.A(_01235_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(net417),
    .A1(net339),
    .S(_01234_),
    .X(_01236_));
 sky130_fd_sc_hd__clkbuf_1 _07528_ (.A(_01236_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _07529_ (.A0(net434),
    .A1(net215),
    .S(_01234_),
    .X(_01237_));
 sky130_fd_sc_hd__clkbuf_1 _07530_ (.A(_01237_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _07531_ (.A0(net73),
    .A1(net348),
    .S(_01234_),
    .X(_01238_));
 sky130_fd_sc_hd__clkbuf_1 _07532_ (.A(net349),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _07533_ (.A0(net384),
    .A1(net334),
    .S(_01234_),
    .X(_01239_));
 sky130_fd_sc_hd__clkbuf_1 _07534_ (.A(_01239_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _07535_ (.A0(net381),
    .A1(net346),
    .S(_01234_),
    .X(_01240_));
 sky130_fd_sc_hd__clkbuf_1 _07536_ (.A(_01240_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _07537_ (.A0(net372),
    .A1(net322),
    .S(_01234_),
    .X(_01241_));
 sky130_fd_sc_hd__clkbuf_1 _07538_ (.A(_01241_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _07539_ (.A0(net375),
    .A1(net236),
    .S(_01234_),
    .X(_01242_));
 sky130_fd_sc_hd__clkbuf_1 _07540_ (.A(_01242_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _07541_ (.A0(net366),
    .A1(net320),
    .S(_01234_),
    .X(_01243_));
 sky130_fd_sc_hd__clkbuf_1 _07542_ (.A(_01243_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _07543_ (.A0(net407),
    .A1(net317),
    .S(_01234_),
    .X(_01244_));
 sky130_fd_sc_hd__clkbuf_1 _07544_ (.A(_01244_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _07545_ (.A0(net415),
    .A1(net278),
    .S(_01012_),
    .X(_01245_));
 sky130_fd_sc_hd__clkbuf_1 _07546_ (.A(_01245_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _07547_ (.A0(net430),
    .A1(net293),
    .S(_01012_),
    .X(_01246_));
 sky130_fd_sc_hd__clkbuf_1 _07548_ (.A(_01246_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _07549_ (.A0(net65),
    .A1(net432),
    .S(_01012_),
    .X(_01247_));
 sky130_fd_sc_hd__clkbuf_1 _07550_ (.A(net433),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _07551_ (.A0(net66),
    .A1(net412),
    .S(_01012_),
    .X(_01248_));
 sky130_fd_sc_hd__clkbuf_1 _07552_ (.A(net413),
    .X(_00067_));
 sky130_fd_sc_hd__clkbuf_4 _07553_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_01249_));
 sky130_fd_sc_hd__buf_4 _07554_ (.A(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__buf_2 _07555_ (.A(net1),
    .X(_01251_));
 sky130_fd_sc_hd__buf_4 _07556_ (.A(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__buf_4 _07557_ (.A(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__and2_1 _07558_ (.A(_01250_),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__clkbuf_1 _07559_ (.A(_01254_),
    .X(_00068_));
 sky130_fd_sc_hd__clkbuf_4 _07560_ (.A(diff_valid),
    .X(_01255_));
 sky130_fd_sc_hd__clkbuf_1 _07561_ (.A(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__clkbuf_1 _07562_ (.A(_01256_),
    .X(_00069_));
 sky130_fd_sc_hd__inv_2 _07563_ (.A(\diff3[17] ),
    .Y(_01257_));
 sky130_fd_sc_hd__a21oi_4 _07564_ (.A1(_01257_),
    .A2(\diff2[17] ),
    .B1(\diff1[17] ),
    .Y(_01258_));
 sky130_fd_sc_hd__o21ai_2 _07565_ (.A1(_01257_),
    .A2(\diff2[17] ),
    .B1(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__inv_2 _07566_ (.A(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__mux2_1 _07567_ (.A0(net206),
    .A1(_01260_),
    .S(_01255_),
    .X(_01261_));
 sky130_fd_sc_hd__clkbuf_1 _07568_ (.A(_01261_),
    .X(_00070_));
 sky130_fd_sc_hd__nor2_1 _07569_ (.A(\diff2[17] ),
    .B(\diff1[17] ),
    .Y(_01262_));
 sky130_fd_sc_hd__mux2_1 _07570_ (.A0(net242),
    .A1(_01262_),
    .S(_01255_),
    .X(_01263_));
 sky130_fd_sc_hd__clkbuf_1 _07571_ (.A(_01263_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(net250),
    .A1(net450),
    .S(_01255_),
    .X(_01264_));
 sky130_fd_sc_hd__clkbuf_1 _07573_ (.A(_01264_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _07574_ (.A0(net292),
    .A1(net360),
    .S(_01255_),
    .X(_01265_));
 sky130_fd_sc_hd__clkbuf_1 _07575_ (.A(_01265_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _07576_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ),
    .A1(net380),
    .S(_01255_),
    .X(_01266_));
 sky130_fd_sc_hd__clkbuf_1 _07577_ (.A(_01266_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _07578_ (.A0(\diff1[3] ),
    .A1(\diff2[3] ),
    .S(_01259_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _07579_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ),
    .A1(_01267_),
    .S(_01255_),
    .X(_01268_));
 sky130_fd_sc_hd__clkbuf_1 _07580_ (.A(_01268_),
    .X(_00075_));
 sky130_fd_sc_hd__and2_1 _07581_ (.A(_01259_),
    .B(_01262_),
    .X(_01269_));
 sky130_fd_sc_hd__clkbuf_4 _07582_ (.A(_01269_),
    .X(_01270_));
 sky130_fd_sc_hd__nor2_1 _07583_ (.A(\diff2[17] ),
    .B(_01259_),
    .Y(_01271_));
 sky130_fd_sc_hd__clkbuf_4 _07584_ (.A(_01271_),
    .X(_01272_));
 sky130_fd_sc_hd__buf_2 _07585_ (.A(\diff2[17] ),
    .X(_01273_));
 sky130_fd_sc_hd__and2_1 _07586_ (.A(_01273_),
    .B(\diff1[4] ),
    .X(_01274_));
 sky130_fd_sc_hd__a221o_1 _07587_ (.A1(\diff2[4] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[4] ),
    .C1(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__clkbuf_4 _07588_ (.A(_01258_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _07589_ (.A0(\r_i_alpha1[4] ),
    .A1(_01275_),
    .S(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _07590_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ),
    .A1(_01277_),
    .S(_01255_),
    .X(_01278_));
 sky130_fd_sc_hd__clkbuf_1 _07591_ (.A(_01278_),
    .X(_00076_));
 sky130_fd_sc_hd__and2_1 _07592_ (.A(_01273_),
    .B(\diff1[5] ),
    .X(_01279_));
 sky130_fd_sc_hd__a221o_1 _07593_ (.A1(\diff2[5] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[5] ),
    .C1(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _07594_ (.A0(\r_i_alpha1[5] ),
    .A1(_01280_),
    .S(_01276_),
    .X(_01281_));
 sky130_fd_sc_hd__clkbuf_4 _07595_ (.A(diff_valid),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _07596_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ),
    .A1(_01281_),
    .S(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__clkbuf_1 _07597_ (.A(_01283_),
    .X(_00077_));
 sky130_fd_sc_hd__and2_1 _07598_ (.A(_01273_),
    .B(\diff1[6] ),
    .X(_01284_));
 sky130_fd_sc_hd__a221o_1 _07599_ (.A1(\diff2[6] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[6] ),
    .C1(_01284_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _07600_ (.A0(\r_i_alpha1[6] ),
    .A1(_01285_),
    .S(_01276_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _07601_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .A1(_01286_),
    .S(_01282_),
    .X(_01287_));
 sky130_fd_sc_hd__clkbuf_1 _07602_ (.A(_01287_),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _07603_ (.A(_01273_),
    .B(\diff1[7] ),
    .X(_01288_));
 sky130_fd_sc_hd__a221o_1 _07604_ (.A1(\diff2[7] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[7] ),
    .C1(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _07605_ (.A0(\r_i_alpha1[7] ),
    .A1(_01289_),
    .S(_01276_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _07606_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ),
    .A1(_01290_),
    .S(_01282_),
    .X(_01291_));
 sky130_fd_sc_hd__clkbuf_1 _07607_ (.A(_01291_),
    .X(_00079_));
 sky130_fd_sc_hd__and2_1 _07608_ (.A(_01273_),
    .B(\diff1[8] ),
    .X(_01292_));
 sky130_fd_sc_hd__a221o_1 _07609_ (.A1(\diff2[8] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[8] ),
    .C1(_01292_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _07610_ (.A0(\r_i_alpha1[8] ),
    .A1(_01293_),
    .S(_01276_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _07611_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ),
    .A1(_01294_),
    .S(_01282_),
    .X(_01295_));
 sky130_fd_sc_hd__clkbuf_1 _07612_ (.A(_01295_),
    .X(_00080_));
 sky130_fd_sc_hd__and2_1 _07613_ (.A(_01273_),
    .B(\diff1[9] ),
    .X(_01296_));
 sky130_fd_sc_hd__a221o_1 _07614_ (.A1(\diff2[9] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[9] ),
    .C1(_01296_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _07615_ (.A0(\r_i_alpha1[9] ),
    .A1(_01297_),
    .S(_01276_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _07616_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ),
    .A1(_01298_),
    .S(_01282_),
    .X(_01299_));
 sky130_fd_sc_hd__clkbuf_1 _07617_ (.A(_01299_),
    .X(_00081_));
 sky130_fd_sc_hd__and2_1 _07618_ (.A(_01273_),
    .B(\diff1[10] ),
    .X(_01300_));
 sky130_fd_sc_hd__a221o_1 _07619_ (.A1(\diff2[10] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[10] ),
    .C1(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _07620_ (.A0(\r_i_alpha1[10] ),
    .A1(_01301_),
    .S(_01276_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _07621_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ),
    .A1(_01302_),
    .S(_01282_),
    .X(_01303_));
 sky130_fd_sc_hd__clkbuf_1 _07622_ (.A(_01303_),
    .X(_00082_));
 sky130_fd_sc_hd__and2_1 _07623_ (.A(_01273_),
    .B(\diff1[11] ),
    .X(_01304_));
 sky130_fd_sc_hd__a221o_1 _07624_ (.A1(\diff2[11] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[11] ),
    .C1(_01304_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _07625_ (.A0(\r_i_alpha1[11] ),
    .A1(_01305_),
    .S(_01276_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _07626_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ),
    .A1(_01306_),
    .S(_01282_),
    .X(_01307_));
 sky130_fd_sc_hd__clkbuf_1 _07627_ (.A(_01307_),
    .X(_00083_));
 sky130_fd_sc_hd__and2_1 _07628_ (.A(_01273_),
    .B(\diff1[12] ),
    .X(_01308_));
 sky130_fd_sc_hd__a221o_1 _07629_ (.A1(\diff2[12] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[12] ),
    .C1(_01308_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _07630_ (.A0(\r_i_alpha1[12] ),
    .A1(_01309_),
    .S(_01276_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _07631_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .A1(_01310_),
    .S(_01282_),
    .X(_01311_));
 sky130_fd_sc_hd__clkbuf_1 _07632_ (.A(_01311_),
    .X(_00084_));
 sky130_fd_sc_hd__and2_1 _07633_ (.A(\diff2[17] ),
    .B(\diff1[13] ),
    .X(_01312_));
 sky130_fd_sc_hd__a221o_1 _07634_ (.A1(\diff2[13] ),
    .A2(_01270_),
    .B1(_01272_),
    .B2(\diff3[13] ),
    .C1(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(\r_i_alpha1[13] ),
    .A1(_01313_),
    .S(_01258_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _07636_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ),
    .A1(_01314_),
    .S(_01282_),
    .X(_01315_));
 sky130_fd_sc_hd__clkbuf_1 _07637_ (.A(_01315_),
    .X(_00085_));
 sky130_fd_sc_hd__and2_1 _07638_ (.A(\diff2[17] ),
    .B(\diff1[14] ),
    .X(_01316_));
 sky130_fd_sc_hd__a221o_1 _07639_ (.A1(\diff2[14] ),
    .A2(_01269_),
    .B1(_01271_),
    .B2(\diff3[14] ),
    .C1(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _07640_ (.A0(\r_i_alpha1[14] ),
    .A1(_01317_),
    .S(_01258_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ),
    .A1(_01318_),
    .S(_01282_),
    .X(_01319_));
 sky130_fd_sc_hd__clkbuf_1 _07642_ (.A(_01319_),
    .X(_00086_));
 sky130_fd_sc_hd__and2_1 _07643_ (.A(\diff2[17] ),
    .B(\diff1[15] ),
    .X(_01320_));
 sky130_fd_sc_hd__a221o_1 _07644_ (.A1(\diff2[15] ),
    .A2(_01269_),
    .B1(_01271_),
    .B2(\diff3[15] ),
    .C1(_01320_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _07645_ (.A0(\r_i_alpha1[15] ),
    .A1(_01321_),
    .S(_01258_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _07646_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ),
    .A1(_01322_),
    .S(diff_valid),
    .X(_01323_));
 sky130_fd_sc_hd__clkbuf_1 _07647_ (.A(_01323_),
    .X(_00087_));
 sky130_fd_sc_hd__and2_1 _07648_ (.A(\diff2[17] ),
    .B(\diff1[16] ),
    .X(_01324_));
 sky130_fd_sc_hd__a221o_1 _07649_ (.A1(\diff2[16] ),
    .A2(_01269_),
    .B1(_01271_),
    .B2(\diff3[16] ),
    .C1(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _07650_ (.A0(\r_i_alpha1[16] ),
    .A1(_01325_),
    .S(_01258_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _07651_ (.A0(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[16] ),
    .A1(_01326_),
    .S(diff_valid),
    .X(_01327_));
 sky130_fd_sc_hd__clkbuf_1 _07652_ (.A(_01327_),
    .X(_00088_));
 sky130_fd_sc_hd__inv_2 _07653_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .Y(_01328_));
 sky130_fd_sc_hd__buf_4 _07654_ (.A(_01328_),
    .X(_01329_));
 sky130_fd_sc_hd__buf_4 _07655_ (.A(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(net178),
    .B(_01255_),
    .Y(_01331_));
 sky130_fd_sc_hd__o22ai_1 _07657_ (.A1(_01330_),
    .A2(_01255_),
    .B1(_01276_),
    .B2(_01331_),
    .Y(_00089_));
 sky130_fd_sc_hd__clkbuf_1 _07658_ (.A(_01059_),
    .X(_01332_));
 sky130_fd_sc_hd__clkbuf_1 _07659_ (.A(_01332_),
    .X(_00090_));
 sky130_fd_sc_hd__clkbuf_4 _07660_ (.A(_00993_),
    .X(_01333_));
 sky130_fd_sc_hd__clkbuf_4 _07661_ (.A(net14),
    .X(_01334_));
 sky130_fd_sc_hd__o21ai_1 _07662_ (.A1(_00991_),
    .A2(_01334_),
    .B1(_00992_),
    .Y(_01335_));
 sky130_fd_sc_hd__a21oi_1 _07663_ (.A1(_00991_),
    .A2(_01334_),
    .B1(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__o21ba_1 _07664_ (.A1(net202),
    .A2(_01333_),
    .B1_N(_01336_),
    .X(_00091_));
 sky130_fd_sc_hd__o21a_1 _07665_ (.A1(_00991_),
    .A2(_01334_),
    .B1(net16),
    .X(_01337_));
 sky130_fd_sc_hd__clkbuf_4 _07666_ (.A(_00992_),
    .X(_01338_));
 sky130_fd_sc_hd__or3_1 _07667_ (.A(_00991_),
    .B(_01334_),
    .C(net16),
    .X(_01339_));
 sky130_fd_sc_hd__nand2_1 _07668_ (.A(_01338_),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__o22a_1 _07669_ (.A1(net228),
    .A2(_01333_),
    .B1(_01337_),
    .B2(_01340_),
    .X(_00092_));
 sky130_fd_sc_hd__or3_2 _07670_ (.A(net15),
    .B(net16),
    .C(net17),
    .X(_01341_));
 sky130_fd_sc_hd__a2bb2o_1 _07671_ (.A1_N(_01334_),
    .A2_N(_01341_),
    .B1(_01339_),
    .B2(net17),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _07672_ (.A0(net347),
    .A1(_01342_),
    .S(_01000_),
    .X(_01343_));
 sky130_fd_sc_hd__clkbuf_1 _07673_ (.A(_01343_),
    .X(_00093_));
 sky130_fd_sc_hd__clkinv_4 _07674_ (.A(_00992_),
    .Y(_01344_));
 sky130_fd_sc_hd__clkbuf_4 _07675_ (.A(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__or3_1 _07676_ (.A(_01334_),
    .B(net18),
    .C(_01341_),
    .X(_01346_));
 sky130_fd_sc_hd__o21a_1 _07677_ (.A1(_01334_),
    .A2(_01341_),
    .B1(net18),
    .X(_01347_));
 sky130_fd_sc_hd__nor2_1 _07678_ (.A(_01344_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__a22o_1 _07679_ (.A1(net190),
    .A2(_01345_),
    .B1(_01346_),
    .B2(_01348_),
    .X(_00094_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(net19),
    .B(_01347_),
    .Y(_01349_));
 sky130_fd_sc_hd__or2_1 _07681_ (.A(net19),
    .B(_01347_),
    .X(_01350_));
 sky130_fd_sc_hd__nand2_1 _07682_ (.A(_01349_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__mux2_1 _07683_ (.A0(net326),
    .A1(_01351_),
    .S(_01000_),
    .X(_01352_));
 sky130_fd_sc_hd__clkbuf_1 _07684_ (.A(_01352_),
    .X(_00095_));
 sky130_fd_sc_hd__or2_1 _07685_ (.A(net20),
    .B(_01350_),
    .X(_01353_));
 sky130_fd_sc_hd__a21oi_1 _07686_ (.A1(net20),
    .A2(_01350_),
    .B1(_01345_),
    .Y(_01354_));
 sky130_fd_sc_hd__o2bb2a_1 _07687_ (.A1_N(_01353_),
    .A2_N(_01354_),
    .B1(net227),
    .B2(_01333_),
    .X(_00096_));
 sky130_fd_sc_hd__and2_1 _07688_ (.A(net4),
    .B(_01353_),
    .X(_01355_));
 sky130_fd_sc_hd__o21ai_1 _07689_ (.A1(net4),
    .A2(_01353_),
    .B1(_01338_),
    .Y(_01356_));
 sky130_fd_sc_hd__a2bb2o_1 _07690_ (.A1_N(_01355_),
    .A2_N(_01356_),
    .B1(net181),
    .B2(_01345_),
    .X(_00097_));
 sky130_fd_sc_hd__xnor2_1 _07691_ (.A(net5),
    .B(_01355_),
    .Y(_01357_));
 sky130_fd_sc_hd__buf_4 _07692_ (.A(_00992_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _07693_ (.A0(net337),
    .A1(_01357_),
    .S(_01358_),
    .X(_01359_));
 sky130_fd_sc_hd__clkbuf_1 _07694_ (.A(_01359_),
    .X(_00098_));
 sky130_fd_sc_hd__o21ai_1 _07695_ (.A1(net5),
    .A2(_01355_),
    .B1(_01003_),
    .Y(_01360_));
 sky130_fd_sc_hd__or3_2 _07696_ (.A(net5),
    .B(_01003_),
    .C(_01355_),
    .X(_01361_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(_01360_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__mux2_1 _07698_ (.A0(net340),
    .A1(_01362_),
    .S(_01358_),
    .X(_01363_));
 sky130_fd_sc_hd__clkbuf_1 _07699_ (.A(_01363_),
    .X(_00099_));
 sky130_fd_sc_hd__xor2_1 _07700_ (.A(net7),
    .B(_01361_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _07701_ (.A0(net345),
    .A1(_01364_),
    .S(_01358_),
    .X(_01365_));
 sky130_fd_sc_hd__clkbuf_1 _07702_ (.A(_01365_),
    .X(_00100_));
 sky130_fd_sc_hd__and3_1 _07703_ (.A(net7),
    .B(net8),
    .C(_01361_),
    .X(_01366_));
 sky130_fd_sc_hd__a21o_1 _07704_ (.A1(net7),
    .A2(_01361_),
    .B1(net8),
    .X(_01367_));
 sky130_fd_sc_hd__nand2_1 _07705_ (.A(_01338_),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__a2bb2o_1 _07706_ (.A1_N(_01366_),
    .A2_N(_01368_),
    .B1(net188),
    .B2(_01345_),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _07707_ (.A(net9),
    .B(_01366_),
    .Y(_01369_));
 sky130_fd_sc_hd__mux2_1 _07708_ (.A0(net362),
    .A1(_01369_),
    .S(_01358_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_1 _07709_ (.A(_01370_),
    .X(_00102_));
 sky130_fd_sc_hd__or3_1 _07710_ (.A(net9),
    .B(net10),
    .C(_01366_),
    .X(_01371_));
 sky130_fd_sc_hd__o21ai_1 _07711_ (.A1(net9),
    .A2(_01366_),
    .B1(net10),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _07712_ (.A(_01371_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__mux2_1 _07713_ (.A0(net392),
    .A1(_01373_),
    .S(_01358_),
    .X(_01374_));
 sky130_fd_sc_hd__clkbuf_1 _07714_ (.A(_01374_),
    .X(_00103_));
 sky130_fd_sc_hd__nor2_1 _07715_ (.A(net11),
    .B(_01371_),
    .Y(_01375_));
 sky130_fd_sc_hd__a21o_1 _07716_ (.A1(net11),
    .A2(_01371_),
    .B1(_01344_),
    .X(_01376_));
 sky130_fd_sc_hd__o22a_1 _07717_ (.A1(net466),
    .A2(_01333_),
    .B1(_01375_),
    .B2(_01376_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _07718_ (.A0(net397),
    .A1(_01334_),
    .S(_01358_),
    .X(_01377_));
 sky130_fd_sc_hd__clkbuf_1 _07719_ (.A(_01377_),
    .X(_00105_));
 sky130_fd_sc_hd__inv_2 _07720_ (.A(_00991_),
    .Y(_01378_));
 sky130_fd_sc_hd__mux2_1 _07721_ (.A0(_01378_),
    .A1(net445),
    .S(_01344_),
    .X(_01379_));
 sky130_fd_sc_hd__clkbuf_1 _07722_ (.A(_01379_),
    .X(_00106_));
 sky130_fd_sc_hd__and2_1 _07723_ (.A(_00991_),
    .B(net16),
    .X(_01380_));
 sky130_fd_sc_hd__o21ai_1 _07724_ (.A1(_00991_),
    .A2(net16),
    .B1(_00993_),
    .Y(_01381_));
 sky130_fd_sc_hd__o22a_1 _07725_ (.A1(net196),
    .A2(_01333_),
    .B1(_01380_),
    .B2(_01381_),
    .X(_00107_));
 sky130_fd_sc_hd__o21a_1 _07726_ (.A1(_00991_),
    .A2(net16),
    .B1(net17),
    .X(_01382_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(_01338_),
    .B(_01341_),
    .Y(_01383_));
 sky130_fd_sc_hd__o22a_1 _07728_ (.A1(net224),
    .A2(_01333_),
    .B1(_01382_),
    .B2(_01383_),
    .X(_00108_));
 sky130_fd_sc_hd__nand2_1 _07729_ (.A(net18),
    .B(_01341_),
    .Y(_01384_));
 sky130_fd_sc_hd__or2_1 _07730_ (.A(net18),
    .B(_01341_),
    .X(_01385_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_01384_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__mux2_1 _07732_ (.A0(net379),
    .A1(_01386_),
    .S(_01358_),
    .X(_01387_));
 sky130_fd_sc_hd__clkbuf_1 _07733_ (.A(_01387_),
    .X(_00109_));
 sky130_fd_sc_hd__or2_1 _07734_ (.A(net19),
    .B(_01385_),
    .X(_01388_));
 sky130_fd_sc_hd__a21oi_1 _07735_ (.A1(net19),
    .A2(_01385_),
    .B1(_01344_),
    .Y(_01389_));
 sky130_fd_sc_hd__a22o_1 _07736_ (.A1(net199),
    .A2(_01345_),
    .B1(_01388_),
    .B2(_01389_),
    .X(_00110_));
 sky130_fd_sc_hd__and3_1 _07737_ (.A(net19),
    .B(net20),
    .C(_01385_),
    .X(_01390_));
 sky130_fd_sc_hd__a21o_1 _07738_ (.A1(net19),
    .A2(_01385_),
    .B1(net20),
    .X(_01391_));
 sky130_fd_sc_hd__nand2_1 _07739_ (.A(_01338_),
    .B(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__o22a_1 _07740_ (.A1(net195),
    .A2(_01338_),
    .B1(_01390_),
    .B2(_01392_),
    .X(_00111_));
 sky130_fd_sc_hd__or2_1 _07741_ (.A(net4),
    .B(_01391_),
    .X(_01393_));
 sky130_fd_sc_hd__a21oi_1 _07742_ (.A1(net4),
    .A2(_01391_),
    .B1(_01344_),
    .Y(_01394_));
 sky130_fd_sc_hd__o2bb2a_1 _07743_ (.A1_N(_01393_),
    .A2_N(_01394_),
    .B1(net239),
    .B2(_01333_),
    .X(_00112_));
 sky130_fd_sc_hd__and2_1 _07744_ (.A(net5),
    .B(_01393_),
    .X(_01395_));
 sky130_fd_sc_hd__o21ai_1 _07745_ (.A1(net5),
    .A2(_01393_),
    .B1(_01338_),
    .Y(_01396_));
 sky130_fd_sc_hd__a2bb2o_1 _07746_ (.A1_N(_01395_),
    .A2_N(_01396_),
    .B1(net194),
    .B2(_01345_),
    .X(_00113_));
 sky130_fd_sc_hd__xnor2_1 _07747_ (.A(_01003_),
    .B(_01395_),
    .Y(_01397_));
 sky130_fd_sc_hd__mux2_1 _07748_ (.A0(net394),
    .A1(_01397_),
    .S(_01358_),
    .X(_01398_));
 sky130_fd_sc_hd__clkbuf_1 _07749_ (.A(_01398_),
    .X(_00114_));
 sky130_fd_sc_hd__o21ai_1 _07750_ (.A1(_01003_),
    .A2(_01395_),
    .B1(net7),
    .Y(_01399_));
 sky130_fd_sc_hd__or3_2 _07751_ (.A(_01003_),
    .B(net7),
    .C(_01395_),
    .X(_01400_));
 sky130_fd_sc_hd__nand2_1 _07752_ (.A(_01399_),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__mux2_1 _07753_ (.A0(net418),
    .A1(_01401_),
    .S(_01358_),
    .X(_01402_));
 sky130_fd_sc_hd__clkbuf_1 _07754_ (.A(_01402_),
    .X(_00115_));
 sky130_fd_sc_hd__xor2_1 _07755_ (.A(net8),
    .B(_01400_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _07756_ (.A0(net472),
    .A1(_01403_),
    .S(_01358_),
    .X(_01404_));
 sky130_fd_sc_hd__clkbuf_1 _07757_ (.A(_01404_),
    .X(_00116_));
 sky130_fd_sc_hd__and3_1 _07758_ (.A(net8),
    .B(net9),
    .C(_01400_),
    .X(_01405_));
 sky130_fd_sc_hd__a21o_1 _07759_ (.A1(net8),
    .A2(_01400_),
    .B1(net9),
    .X(_01406_));
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(_01338_),
    .B(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__a2bb2o_1 _07761_ (.A1_N(_01405_),
    .A2_N(_01407_),
    .B1(net262),
    .B2(_01345_),
    .X(_00117_));
 sky130_fd_sc_hd__or2_1 _07762_ (.A(net10),
    .B(_01405_),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _07763_ (.A(net10),
    .B(_01405_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_1 _07764_ (.A(_01408_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__buf_4 _07765_ (.A(_00992_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _07766_ (.A0(net438),
    .A1(_01410_),
    .S(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__clkbuf_1 _07767_ (.A(_01412_),
    .X(_00118_));
 sky130_fd_sc_hd__xnor2_1 _07768_ (.A(net11),
    .B(_01408_),
    .Y(_01413_));
 sky130_fd_sc_hd__mux2_1 _07769_ (.A0(_01273_),
    .A1(_01413_),
    .S(_01411_),
    .X(_01414_));
 sky130_fd_sc_hd__clkbuf_1 _07770_ (.A(_01414_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _07771_ (.A0(net450),
    .A1(net3),
    .S(_01411_),
    .X(_01415_));
 sky130_fd_sc_hd__clkbuf_1 _07772_ (.A(_01415_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _07773_ (.A0(net360),
    .A1(net12),
    .S(_01411_),
    .X(_01416_));
 sky130_fd_sc_hd__clkbuf_1 _07774_ (.A(_01416_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _07775_ (.A0(net380),
    .A1(net13),
    .S(_01411_),
    .X(_01417_));
 sky130_fd_sc_hd__clkbuf_1 _07776_ (.A(_01417_),
    .X(_00122_));
 sky130_fd_sc_hd__inv_2 _07777_ (.A(_01334_),
    .Y(_01418_));
 sky130_fd_sc_hd__mux2_1 _07778_ (.A0(_01418_),
    .A1(net404),
    .S(_01344_),
    .X(_01419_));
 sky130_fd_sc_hd__clkbuf_1 _07779_ (.A(_01419_),
    .X(_00123_));
 sky130_fd_sc_hd__a21o_1 _07780_ (.A1(net189),
    .A2(_01345_),
    .B1(_01336_),
    .X(_00124_));
 sky130_fd_sc_hd__and3_1 _07781_ (.A(_00991_),
    .B(_01334_),
    .C(net16),
    .X(_01420_));
 sky130_fd_sc_hd__a21o_1 _07782_ (.A1(net15),
    .A2(net14),
    .B1(net16),
    .X(_01421_));
 sky130_fd_sc_hd__nand2_1 _07783_ (.A(_01338_),
    .B(_01421_),
    .Y(_01422_));
 sky130_fd_sc_hd__o22a_1 _07784_ (.A1(net232),
    .A2(_01338_),
    .B1(_01420_),
    .B2(_01422_),
    .X(_00125_));
 sky130_fd_sc_hd__or2_1 _07785_ (.A(net17),
    .B(_01421_),
    .X(_01423_));
 sky130_fd_sc_hd__a21oi_1 _07786_ (.A1(net17),
    .A2(_01421_),
    .B1(_01344_),
    .Y(_01424_));
 sky130_fd_sc_hd__o2bb2a_1 _07787_ (.A1_N(_01423_),
    .A2_N(_01424_),
    .B1(net247),
    .B2(_01333_),
    .X(_00126_));
 sky130_fd_sc_hd__xor2_1 _07788_ (.A(net18),
    .B(_01423_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _07789_ (.A0(net425),
    .A1(_01425_),
    .S(_01411_),
    .X(_01426_));
 sky130_fd_sc_hd__clkbuf_1 _07790_ (.A(_01426_),
    .X(_00127_));
 sky130_fd_sc_hd__a21oi_1 _07791_ (.A1(net18),
    .A2(_01423_),
    .B1(net19),
    .Y(_01427_));
 sky130_fd_sc_hd__and3_1 _07792_ (.A(net18),
    .B(net19),
    .C(_01423_),
    .X(_01428_));
 sky130_fd_sc_hd__nor2_1 _07793_ (.A(_01427_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__mux2_1 _07794_ (.A0(net390),
    .A1(_01429_),
    .S(_01411_),
    .X(_01430_));
 sky130_fd_sc_hd__clkbuf_1 _07795_ (.A(_01430_),
    .X(_00128_));
 sky130_fd_sc_hd__or2_2 _07796_ (.A(net20),
    .B(_01428_),
    .X(_01431_));
 sky130_fd_sc_hd__a21oi_1 _07797_ (.A1(net20),
    .A2(_01428_),
    .B1(_01344_),
    .Y(_01432_));
 sky130_fd_sc_hd__o2bb2a_1 _07798_ (.A1_N(_01431_),
    .A2_N(_01432_),
    .B1(net248),
    .B2(_01333_),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(net4),
    .B(_01431_),
    .Y(_01433_));
 sky130_fd_sc_hd__o21a_1 _07800_ (.A1(net4),
    .A2(_01431_),
    .B1(_00993_),
    .X(_01434_));
 sky130_fd_sc_hd__a22o_1 _07801_ (.A1(net198),
    .A2(_01345_),
    .B1(_01433_),
    .B2(_01434_),
    .X(_00130_));
 sky130_fd_sc_hd__and3_2 _07802_ (.A(net4),
    .B(net5),
    .C(_01431_),
    .X(_01435_));
 sky130_fd_sc_hd__a21oi_1 _07803_ (.A1(net4),
    .A2(_01431_),
    .B1(net5),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_1 _07804_ (.A(_01435_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__mux2_1 _07805_ (.A0(net382),
    .A1(_01437_),
    .S(_01411_),
    .X(_01438_));
 sky130_fd_sc_hd__clkbuf_1 _07806_ (.A(_01438_),
    .X(_00131_));
 sky130_fd_sc_hd__xnor2_1 _07807_ (.A(_01003_),
    .B(_01435_),
    .Y(_01439_));
 sky130_fd_sc_hd__mux2_1 _07808_ (.A0(net383),
    .A1(_01439_),
    .S(_01411_),
    .X(_01440_));
 sky130_fd_sc_hd__clkbuf_1 _07809_ (.A(_01440_),
    .X(_00132_));
 sky130_fd_sc_hd__o21ai_2 _07810_ (.A1(_01003_),
    .A2(_01435_),
    .B1(net7),
    .Y(_01441_));
 sky130_fd_sc_hd__o31a_1 _07811_ (.A1(_01003_),
    .A2(net7),
    .A3(_01435_),
    .B1(_00993_),
    .X(_01442_));
 sky130_fd_sc_hd__a22o_1 _07812_ (.A1(net200),
    .A2(_01345_),
    .B1(_01441_),
    .B2(_01442_),
    .X(_00133_));
 sky130_fd_sc_hd__xor2_1 _07813_ (.A(net8),
    .B(_01441_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _07814_ (.A0(net426),
    .A1(_01443_),
    .S(_01411_),
    .X(_01444_));
 sky130_fd_sc_hd__clkbuf_1 _07815_ (.A(_01444_),
    .X(_00134_));
 sky130_fd_sc_hd__or2b_1 _07816_ (.A(net8),
    .B_N(_01441_),
    .X(_01445_));
 sky130_fd_sc_hd__xnor2_1 _07817_ (.A(net9),
    .B(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__mux2_1 _07818_ (.A0(net396),
    .A1(_01446_),
    .S(_00992_),
    .X(_01447_));
 sky130_fd_sc_hd__clkbuf_1 _07819_ (.A(_01447_),
    .X(_00135_));
 sky130_fd_sc_hd__or3_1 _07820_ (.A(net9),
    .B(net10),
    .C(_01445_),
    .X(_01448_));
 sky130_fd_sc_hd__o21ai_1 _07821_ (.A1(net9),
    .A2(_01445_),
    .B1(net10),
    .Y(_01449_));
 sky130_fd_sc_hd__and2_1 _07822_ (.A(net361),
    .B(_01344_),
    .X(_01450_));
 sky130_fd_sc_hd__a31o_1 _07823_ (.A1(_01333_),
    .A2(_01448_),
    .A3(_01449_),
    .B1(_01450_),
    .X(_00136_));
 sky130_fd_sc_hd__xor2_1 _07824_ (.A(net11),
    .B(_01449_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _07825_ (.A0(net502),
    .A1(_01451_),
    .S(_00992_),
    .X(_01452_));
 sky130_fd_sc_hd__clkbuf_1 _07826_ (.A(_01452_),
    .X(_00137_));
 sky130_fd_sc_hd__inv_2 _07827_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ),
    .Y(_01453_));
 sky130_fd_sc_hd__clkbuf_4 _07828_ (.A(_01453_),
    .X(_01454_));
 sky130_fd_sc_hd__clkbuf_4 _07829_ (.A(_01251_),
    .X(_01455_));
 sky130_fd_sc_hd__buf_4 _07830_ (.A(_01455_),
    .X(_01456_));
 sky130_fd_sc_hd__clkbuf_4 _07831_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ),
    .X(_01457_));
 sky130_fd_sc_hd__or2_1 _07832_ (.A(net203),
    .B(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__o211a_1 _07833_ (.A1(_01454_),
    .A2(net206),
    .B1(_01456_),
    .C1(_01458_),
    .X(_00138_));
 sky130_fd_sc_hd__or2_1 _07834_ (.A(net159),
    .B(_01457_),
    .X(_01459_));
 sky130_fd_sc_hd__o211a_1 _07835_ (.A1(_01454_),
    .A2(net242),
    .B1(_01456_),
    .C1(_01459_),
    .X(_00139_));
 sky130_fd_sc_hd__clkbuf_4 _07836_ (.A(_01455_),
    .X(_01460_));
 sky130_fd_sc_hd__or2_1 _07837_ (.A(net165),
    .B(_01457_),
    .X(_01461_));
 sky130_fd_sc_hd__o211a_1 _07838_ (.A1(_01454_),
    .A2(net250),
    .B1(_01460_),
    .C1(_01461_),
    .X(_00140_));
 sky130_fd_sc_hd__or2_1 _07839_ (.A(net164),
    .B(_01457_),
    .X(_01462_));
 sky130_fd_sc_hd__o211a_1 _07840_ (.A1(_01454_),
    .A2(net292),
    .B1(_01460_),
    .C1(_01462_),
    .X(_00141_));
 sky130_fd_sc_hd__clkbuf_4 _07841_ (.A(_01457_),
    .X(_01463_));
 sky130_fd_sc_hd__clkbuf_4 _07842_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ),
    .X(_01464_));
 sky130_fd_sc_hd__clkbuf_4 _07843_ (.A(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__nand2_1 _07844_ (.A(_01465_),
    .B(net401),
    .Y(_01466_));
 sky130_fd_sc_hd__o211a_1 _07845_ (.A1(_01463_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .B1(_01460_),
    .C1(_01466_),
    .X(_00142_));
 sky130_fd_sc_hd__clkbuf_4 _07846_ (.A(_01464_),
    .X(_01467_));
 sky130_fd_sc_hd__nand2_1 _07847_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ),
    .Y(_01468_));
 sky130_fd_sc_hd__or2_1 _07848_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ),
    .X(_01469_));
 sky130_fd_sc_hd__clkbuf_4 _07849_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .X(_01470_));
 sky130_fd_sc_hd__a21oi_1 _07850_ (.A1(_01468_),
    .A2(_01469_),
    .B1(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__clkbuf_4 _07851_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .X(_01472_));
 sky130_fd_sc_hd__a31o_1 _07852_ (.A1(_01472_),
    .A2(_01468_),
    .A3(_01469_),
    .B1(_01453_),
    .X(_01473_));
 sky130_fd_sc_hd__clkbuf_8 _07853_ (.A(_01251_),
    .X(_01474_));
 sky130_fd_sc_hd__buf_4 _07854_ (.A(_01474_),
    .X(_01475_));
 sky130_fd_sc_hd__o221a_1 _07855_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ),
    .B1(_01471_),
    .B2(_01473_),
    .C1(_01475_),
    .X(_00143_));
 sky130_fd_sc_hd__and3_1 _07856_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ),
    .C(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ),
    .X(_01476_));
 sky130_fd_sc_hd__a21oi_1 _07857_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ),
    .Y(_01477_));
 sky130_fd_sc_hd__or2_1 _07858_ (.A(_01476_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__nor2_1 _07859_ (.A(_01471_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__clkbuf_4 _07860_ (.A(_01453_),
    .X(_01480_));
 sky130_fd_sc_hd__a21o_1 _07861_ (.A1(_01471_),
    .A2(_01478_),
    .B1(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__o221a_1 _07862_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ),
    .B1(_01479_),
    .B2(_01481_),
    .C1(_01475_),
    .X(_00144_));
 sky130_fd_sc_hd__nand2_1 _07863_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .B(_01476_),
    .Y(_01482_));
 sky130_fd_sc_hd__o31a_1 _07864_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ),
    .A3(_01469_),
    .B1(_01482_),
    .X(_01483_));
 sky130_fd_sc_hd__and2_1 _07865_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__buf_4 _07866_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ),
    .X(_01485_));
 sky130_fd_sc_hd__o21ai_1 _07867_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ),
    .A2(_01483_),
    .B1(_01485_),
    .Y(_01486_));
 sky130_fd_sc_hd__o221a_1 _07868_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ),
    .B1(_01484_),
    .B2(_01486_),
    .C1(_01475_),
    .X(_00145_));
 sky130_fd_sc_hd__and2_1 _07869_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ),
    .B(_01476_),
    .X(_01487_));
 sky130_fd_sc_hd__or2_1 _07870_ (.A(_01328_),
    .B(_01487_),
    .X(_01488_));
 sky130_fd_sc_hd__or3_1 _07871_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ),
    .C(_01469_),
    .X(_01489_));
 sky130_fd_sc_hd__nand2_1 _07872_ (.A(_01328_),
    .B(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__a21oi_1 _07873_ (.A1(_01488_),
    .A2(_01490_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .Y(_01491_));
 sky130_fd_sc_hd__a31o_1 _07874_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .A2(_01488_),
    .A3(_01490_),
    .B1(_01453_),
    .X(_01492_));
 sky130_fd_sc_hd__o221a_1 _07875_ (.A1(_01467_),
    .A2(net528),
    .B1(_01491_),
    .B2(_01492_),
    .C1(_01475_),
    .X(_00146_));
 sky130_fd_sc_hd__inv_2 _07876_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ),
    .Y(_01493_));
 sky130_fd_sc_hd__mux2_1 _07877_ (.A0(_01488_),
    .A1(_01490_),
    .S(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .X(_01494_));
 sky130_fd_sc_hd__o21ai_1 _07878_ (.A1(_01493_),
    .A2(_01494_),
    .B1(_01464_),
    .Y(_01495_));
 sky130_fd_sc_hd__a21o_1 _07879_ (.A1(_01493_),
    .A2(_01494_),
    .B1(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__o211a_1 _07880_ (.A1(_01463_),
    .A2(net546),
    .B1(_01460_),
    .C1(_01496_),
    .X(_00147_));
 sky130_fd_sc_hd__o21ai_1 _07881_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .A2(_01487_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ),
    .Y(_01497_));
 sky130_fd_sc_hd__a21o_1 _07882_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .A2(_01489_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _07883_ (.A0(_01497_),
    .A1(_01498_),
    .S(_01329_),
    .X(_01499_));
 sky130_fd_sc_hd__nor2_1 _07884_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__a21o_1 _07885_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ),
    .A2(_01499_),
    .B1(_01480_),
    .X(_01501_));
 sky130_fd_sc_hd__o221a_1 _07886_ (.A1(_01467_),
    .A2(net629),
    .B1(_01500_),
    .B2(_01501_),
    .C1(_01475_),
    .X(_00148_));
 sky130_fd_sc_hd__o211a_1 _07887_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ),
    .A2(_01487_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ),
    .C1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ),
    .X(_01502_));
 sky130_fd_sc_hd__o21ai_1 _07888_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ),
    .A2(_01498_),
    .B1(_01328_),
    .Y(_01503_));
 sky130_fd_sc_hd__o21a_1 _07889_ (.A1(_01329_),
    .A2(_01502_),
    .B1(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__o21ai_1 _07890_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ),
    .A2(_01504_),
    .B1(_01464_),
    .Y(_01505_));
 sky130_fd_sc_hd__a21o_1 _07891_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ),
    .A2(_01504_),
    .B1(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__o211a_1 _07892_ (.A1(_01463_),
    .A2(net500),
    .B1(_01460_),
    .C1(_01506_),
    .X(_00149_));
 sky130_fd_sc_hd__inv_2 _07893_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ),
    .Y(_01507_));
 sky130_fd_sc_hd__or2_1 _07894_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ),
    .B(_01502_),
    .X(_01508_));
 sky130_fd_sc_hd__a22oi_2 _07895_ (.A1(_01329_),
    .A2(_01507_),
    .B1(_01503_),
    .B2(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _07896_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__a21o_1 _07897_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ),
    .A2(_01509_),
    .B1(_01480_),
    .X(_01511_));
 sky130_fd_sc_hd__buf_6 _07898_ (.A(_01252_),
    .X(_01512_));
 sky130_fd_sc_hd__clkbuf_4 _07899_ (.A(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__o221a_1 _07900_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_01510_),
    .B2(_01511_),
    .C1(_01513_),
    .X(_00150_));
 sky130_fd_sc_hd__o21a_1 _07901_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ),
    .A2(_01498_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ),
    .X(_01514_));
 sky130_fd_sc_hd__or2_1 _07902_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ),
    .B(_01514_),
    .X(_01515_));
 sky130_fd_sc_hd__nand2_1 _07903_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ),
    .B(_01508_),
    .Y(_01516_));
 sky130_fd_sc_hd__mux2_1 _07904_ (.A0(_01515_),
    .A1(_01516_),
    .S(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .X(_01517_));
 sky130_fd_sc_hd__nor2_1 _07905_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21o_1 _07906_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ),
    .A2(_01517_),
    .B1(_01480_),
    .X(_01519_));
 sky130_fd_sc_hd__o221a_1 _07907_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[11] ),
    .B1(_01518_),
    .B2(_01519_),
    .C1(_01513_),
    .X(_00151_));
 sky130_fd_sc_hd__and3_1 _07908_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ),
    .C(_01508_),
    .X(_01520_));
 sky130_fd_sc_hd__or2_1 _07909_ (.A(_01328_),
    .B(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__or2_1 _07910_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ),
    .B(_01515_),
    .X(_01522_));
 sky130_fd_sc_hd__nand2_1 _07911_ (.A(_01328_),
    .B(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__a21oi_1 _07912_ (.A1(_01521_),
    .A2(_01523_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .Y(_01524_));
 sky130_fd_sc_hd__a31o_1 _07913_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .A2(_01521_),
    .A3(_01523_),
    .B1(_01453_),
    .X(_01525_));
 sky130_fd_sc_hd__o221a_1 _07914_ (.A1(_01467_),
    .A2(net559),
    .B1(_01524_),
    .B2(_01525_),
    .C1(_01513_),
    .X(_00152_));
 sky130_fd_sc_hd__and2_1 _07915_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .B(_01523_),
    .X(_01526_));
 sky130_fd_sc_hd__and2b_1 _07916_ (.A_N(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .B(_01521_),
    .X(_01527_));
 sky130_fd_sc_hd__o21a_1 _07917_ (.A1(_01526_),
    .A2(_01527_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ),
    .X(_01528_));
 sky130_fd_sc_hd__buf_4 _07918_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ),
    .X(_01529_));
 sky130_fd_sc_hd__o31ai_1 _07919_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ),
    .A2(_01526_),
    .A3(_01527_),
    .B1(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__o221a_1 _07920_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_01528_),
    .B2(_01530_),
    .C1(_01513_),
    .X(_00153_));
 sky130_fd_sc_hd__and3_1 _07921_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ),
    .C(_01522_),
    .X(_01531_));
 sky130_fd_sc_hd__nor2_1 _07922_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__inv_2 _07923_ (.A(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__or3_1 _07924_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ),
    .C(_01520_),
    .X(_01534_));
 sky130_fd_sc_hd__nand2_1 _07925_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__a21oi_1 _07926_ (.A1(_01533_),
    .A2(_01535_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _07927_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ),
    .B(_01535_),
    .Y(_01537_));
 sky130_fd_sc_hd__o21ai_1 _07928_ (.A1(_01532_),
    .A2(_01537_),
    .B1(_01485_),
    .Y(_01538_));
 sky130_fd_sc_hd__o221a_1 _07929_ (.A1(_01467_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_01536_),
    .B2(_01538_),
    .C1(_01513_),
    .X(_00154_));
 sky130_fd_sc_hd__clkbuf_4 _07930_ (.A(_01464_),
    .X(_01539_));
 sky130_fd_sc_hd__o21ai_1 _07931_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ),
    .A2(_01532_),
    .B1(_01537_),
    .Y(_01540_));
 sky130_fd_sc_hd__and2_1 _07932_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__o21ai_1 _07933_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ),
    .A2(_01540_),
    .B1(_01529_),
    .Y(_01542_));
 sky130_fd_sc_hd__o221a_1 _07934_ (.A1(_01539_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_01541_),
    .B2(_01542_),
    .C1(_01513_),
    .X(_00155_));
 sky130_fd_sc_hd__o31a_1 _07935_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ),
    .A3(_01531_),
    .B1(_01328_),
    .X(_01543_));
 sky130_fd_sc_hd__a31o_1 _07936_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ),
    .A3(_01534_),
    .B1(_01328_),
    .X(_01544_));
 sky130_fd_sc_hd__or2b_1 _07937_ (.A(_01543_),
    .B_N(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__nor2_1 _07938_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[16] ),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__a21o_1 _07939_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[16] ),
    .A2(_01545_),
    .B1(_01480_),
    .X(_01547_));
 sky130_fd_sc_hd__o221a_1 _07940_ (.A1(_01539_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[16] ),
    .B1(_01546_),
    .B2(_01547_),
    .C1(_01513_),
    .X(_00156_));
 sky130_fd_sc_hd__a21oi_1 _07941_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[16] ),
    .A2(_01544_),
    .B1(_01543_),
    .Y(_01548_));
 sky130_fd_sc_hd__buf_2 _07942_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_01549_));
 sky130_fd_sc_hd__buf_2 _07943_ (.A(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__or2_1 _07944_ (.A(_01464_),
    .B(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__buf_4 _07945_ (.A(_01455_),
    .X(_01552_));
 sky130_fd_sc_hd__o211a_1 _07946_ (.A1(_01454_),
    .A2(_01548_),
    .B1(_01551_),
    .C1(_01552_),
    .X(_00157_));
 sky130_fd_sc_hd__and2b_1 _07947_ (.A_N(net21),
    .B(net39),
    .X(_01553_));
 sky130_fd_sc_hd__or2b_1 _07948_ (.A(net39),
    .B_N(net21),
    .X(_01554_));
 sky130_fd_sc_hd__nand2_1 _07949_ (.A(_01485_),
    .B(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__o221a_1 _07950_ (.A1(_01539_),
    .A2(net555),
    .B1(_01553_),
    .B2(_01555_),
    .C1(_01513_),
    .X(_00158_));
 sky130_fd_sc_hd__buf_4 _07951_ (.A(_01470_),
    .X(_01556_));
 sky130_fd_sc_hd__xor2_4 _07952_ (.A(net30),
    .B(net48),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_1 _07953_ (.A(net21),
    .B(net39),
    .Y(_01558_));
 sky130_fd_sc_hd__xor2_2 _07954_ (.A(_01557_),
    .B(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__a21oi_1 _07955_ (.A1(net21),
    .A2(_01556_),
    .B1(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__a31o_1 _07956_ (.A1(net21),
    .A2(_01472_),
    .A3(_01559_),
    .B1(_01453_),
    .X(_01561_));
 sky130_fd_sc_hd__o221a_1 _07957_ (.A1(_01539_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B1(_01560_),
    .B2(_01561_),
    .C1(_01513_),
    .X(_00159_));
 sky130_fd_sc_hd__clkbuf_4 _07958_ (.A(_01472_),
    .X(_01562_));
 sky130_fd_sc_hd__and2b_1 _07959_ (.A_N(net49),
    .B(net31),
    .X(_01563_));
 sky130_fd_sc_hd__and2b_1 _07960_ (.A_N(net31),
    .B(net49),
    .X(_01564_));
 sky130_fd_sc_hd__nor2_2 _07961_ (.A(_01563_),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__and2_1 _07962_ (.A(net30),
    .B(net48),
    .X(_01566_));
 sky130_fd_sc_hd__a31oi_4 _07963_ (.A1(net21),
    .A2(net39),
    .A3(_01557_),
    .B1(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__xnor2_2 _07964_ (.A(_01565_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__or2b_1 _07965_ (.A(net48),
    .B_N(net30),
    .X(_01569_));
 sky130_fd_sc_hd__and2b_1 _07966_ (.A_N(net30),
    .B(net48),
    .X(_01570_));
 sky130_fd_sc_hd__a21o_1 _07967_ (.A1(_01554_),
    .A2(_01569_),
    .B1(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__buf_4 _07968_ (.A(_01328_),
    .X(_01572_));
 sky130_fd_sc_hd__a21oi_1 _07969_ (.A1(_01565_),
    .A2(_01571_),
    .B1(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__o21ai_1 _07970_ (.A1(_01565_),
    .A2(_01571_),
    .B1(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__o211ai_2 _07971_ (.A1(_01562_),
    .A2(_01568_),
    .B1(_01574_),
    .C1(_01485_),
    .Y(_01575_));
 sky130_fd_sc_hd__o211a_1 _07972_ (.A1(_01463_),
    .A2(net459),
    .B1(_01460_),
    .C1(_01575_),
    .X(_00160_));
 sky130_fd_sc_hd__and2b_1 _07973_ (.A_N(net32),
    .B(net50),
    .X(_01576_));
 sky130_fd_sc_hd__or2b_1 _07974_ (.A(net50),
    .B_N(net32),
    .X(_01577_));
 sky130_fd_sc_hd__or2b_1 _07975_ (.A(_01576_),
    .B_N(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__clkbuf_2 _07976_ (.A(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__nand2_1 _07977_ (.A(net31),
    .B(net49),
    .Y(_01580_));
 sky130_fd_sc_hd__o21ai_1 _07978_ (.A1(_01565_),
    .A2(_01567_),
    .B1(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__xnor2_1 _07979_ (.A(_01579_),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _07980_ (.A(_01562_),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__a21o_1 _07981_ (.A1(_01565_),
    .A2(_01571_),
    .B1(_01564_),
    .X(_01584_));
 sky130_fd_sc_hd__xnor2_1 _07982_ (.A(_01579_),
    .B(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__a21o_1 _07983_ (.A1(_01556_),
    .A2(_01585_),
    .B1(_01480_),
    .X(_01586_));
 sky130_fd_sc_hd__o221a_1 _07984_ (.A1(_01539_),
    .A2(net613),
    .B1(_01583_),
    .B2(_01586_),
    .C1(_01513_),
    .X(_00161_));
 sky130_fd_sc_hd__or2b_1 _07985_ (.A(net51),
    .B_N(net33),
    .X(_01587_));
 sky130_fd_sc_hd__or2b_2 _07986_ (.A(net33),
    .B_N(net51),
    .X(_01588_));
 sky130_fd_sc_hd__nand2_4 _07987_ (.A(_01587_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__and2_1 _07988_ (.A(net32),
    .B(net50),
    .X(_01590_));
 sky130_fd_sc_hd__a21o_1 _07989_ (.A1(_01579_),
    .A2(_01581_),
    .B1(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _07990_ (.A(_01589_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__a21oi_2 _07991_ (.A1(_01577_),
    .A2(_01584_),
    .B1(_01576_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _07992_ (.A(_01589_),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__a21o_1 _07993_ (.A1(_01589_),
    .A2(_01593_),
    .B1(_01572_),
    .X(_01595_));
 sky130_fd_sc_hd__o221ai_2 _07994_ (.A1(_01556_),
    .A2(_01592_),
    .B1(_01594_),
    .B2(_01595_),
    .C1(_01485_),
    .Y(_01596_));
 sky130_fd_sc_hd__o211a_1 _07995_ (.A1(_01463_),
    .A2(net638),
    .B1(_01460_),
    .C1(_01596_),
    .X(_00162_));
 sky130_fd_sc_hd__or2b_1 _07996_ (.A(net34),
    .B_N(net52),
    .X(_01597_));
 sky130_fd_sc_hd__or2b_2 _07997_ (.A(net52),
    .B_N(net34),
    .X(_01598_));
 sky130_fd_sc_hd__and2_1 _07998_ (.A(_01597_),
    .B(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__and2_1 _07999_ (.A(net33),
    .B(net51),
    .X(_01600_));
 sky130_fd_sc_hd__a21oi_1 _08000_ (.A1(_01589_),
    .A2(_01591_),
    .B1(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__xnor2_1 _08001_ (.A(_01599_),
    .B(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__nand2_1 _08002_ (.A(_01597_),
    .B(_01598_),
    .Y(_01603_));
 sky130_fd_sc_hd__o21a_1 _08003_ (.A1(_01589_),
    .A2(_01593_),
    .B1(_01588_),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _08004_ (.A(_01603_),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__mux2_1 _08005_ (.A0(_01602_),
    .A1(_01605_),
    .S(_01470_),
    .X(_01606_));
 sky130_fd_sc_hd__nand2_1 _08006_ (.A(_01465_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__o211a_1 _08007_ (.A1(_01463_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ),
    .B1(_01460_),
    .C1(_01607_),
    .X(_00163_));
 sky130_fd_sc_hd__inv_2 _08008_ (.A(net53),
    .Y(_01608_));
 sky130_fd_sc_hd__and2_1 _08009_ (.A(net35),
    .B(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__nor2_1 _08010_ (.A(net35),
    .B(_01608_),
    .Y(_01610_));
 sky130_fd_sc_hd__or2_1 _08011_ (.A(_01609_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__buf_2 _08012_ (.A(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__inv_2 _08013_ (.A(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__inv_2 _08014_ (.A(_01598_),
    .Y(_01614_));
 sky130_fd_sc_hd__o211a_1 _08015_ (.A1(_01589_),
    .A2(_01593_),
    .B1(_01597_),
    .C1(_01588_),
    .X(_01615_));
 sky130_fd_sc_hd__nor2_1 _08016_ (.A(_01614_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__xnor2_1 _08017_ (.A(_01613_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__and2_1 _08018_ (.A(net34),
    .B(net52),
    .X(_01618_));
 sky130_fd_sc_hd__and2_1 _08019_ (.A(_01603_),
    .B(_01600_),
    .X(_01619_));
 sky130_fd_sc_hd__a311o_1 _08020_ (.A1(_01589_),
    .A2(_01591_),
    .A3(_01603_),
    .B1(_01618_),
    .C1(_01619_),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_1 _08021_ (.A(_01612_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__o21a_1 _08022_ (.A1(_01472_),
    .A2(_01621_),
    .B1(_01464_),
    .X(_01622_));
 sky130_fd_sc_hd__o21ai_1 _08023_ (.A1(_01330_),
    .A2(_01617_),
    .B1(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__o211a_1 _08024_ (.A1(_01463_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_01460_),
    .C1(_01623_),
    .X(_00164_));
 sky130_fd_sc_hd__inv_2 _08025_ (.A(net54),
    .Y(_01624_));
 sky130_fd_sc_hd__or2_2 _08026_ (.A(net36),
    .B(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__nand2_1 _08027_ (.A(net36),
    .B(_01624_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_2 _08028_ (.A(_01625_),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__and2_1 _08029_ (.A(net35),
    .B(net53),
    .X(_01628_));
 sky130_fd_sc_hd__a21o_1 _08030_ (.A1(_01612_),
    .A2(_01620_),
    .B1(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__xnor2_1 _08031_ (.A(_01627_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__a21oi_1 _08032_ (.A1(_01613_),
    .A2(_01616_),
    .B1(_01610_),
    .Y(_01631_));
 sky130_fd_sc_hd__xnor2_1 _08033_ (.A(_01627_),
    .B(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__mux2_1 _08034_ (.A0(_01630_),
    .A1(_01632_),
    .S(_01470_),
    .X(_01633_));
 sky130_fd_sc_hd__nand2_1 _08035_ (.A(_01465_),
    .B(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__o211a_1 _08036_ (.A1(_01463_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_01460_),
    .C1(_01634_),
    .X(_00165_));
 sky130_fd_sc_hd__clkbuf_4 _08037_ (.A(_01455_),
    .X(_01635_));
 sky130_fd_sc_hd__or2b_2 _08038_ (.A(net55),
    .B_N(net37),
    .X(_01636_));
 sky130_fd_sc_hd__or2b_2 _08039_ (.A(net37),
    .B_N(net55),
    .X(_01637_));
 sky130_fd_sc_hd__nand2_4 _08040_ (.A(_01636_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__and2_1 _08041_ (.A(net36),
    .B(net54),
    .X(_01639_));
 sky130_fd_sc_hd__a31o_1 _08042_ (.A1(net35),
    .A2(net53),
    .A3(_01627_),
    .B1(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__a31o_2 _08043_ (.A1(_01612_),
    .A2(_01620_),
    .A3(_01627_),
    .B1(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__xnor2_2 _08044_ (.A(_01638_),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor2_1 _08045_ (.A(_01612_),
    .B(_01627_),
    .Y(_01643_));
 sky130_fd_sc_hd__inv_2 _08046_ (.A(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _08047_ (.A(_01610_),
    .B(_01626_),
    .Y(_01645_));
 sky130_fd_sc_hd__o31a_1 _08048_ (.A1(_01614_),
    .A2(_01615_),
    .A3(_01644_),
    .B1(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__and2_1 _08049_ (.A(_01625_),
    .B(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__nor2_1 _08050_ (.A(_01638_),
    .B(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__a31o_1 _08051_ (.A1(_01625_),
    .A2(_01638_),
    .A3(_01646_),
    .B1(_01572_),
    .X(_01649_));
 sky130_fd_sc_hd__o221ai_2 _08052_ (.A1(_01556_),
    .A2(_01642_),
    .B1(_01648_),
    .B2(_01649_),
    .C1(_01485_),
    .Y(_01650_));
 sky130_fd_sc_hd__o211a_1 _08053_ (.A1(_01463_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_01635_),
    .C1(_01650_),
    .X(_00166_));
 sky130_fd_sc_hd__and2b_1 _08054_ (.A_N(net56),
    .B(net38),
    .X(_01651_));
 sky130_fd_sc_hd__and2b_1 _08055_ (.A_N(net38),
    .B(net56),
    .X(_01652_));
 sky130_fd_sc_hd__nor2_1 _08056_ (.A(_01651_),
    .B(_01652_),
    .Y(_01653_));
 sky130_fd_sc_hd__and2_1 _08057_ (.A(net37),
    .B(net55),
    .X(_01654_));
 sky130_fd_sc_hd__a21oi_1 _08058_ (.A1(_01638_),
    .A2(_01641_),
    .B1(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__xnor2_1 _08059_ (.A(_01653_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _08060_ (.A(_01562_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__o21a_1 _08061_ (.A1(_01638_),
    .A2(_01647_),
    .B1(_01637_),
    .X(_01658_));
 sky130_fd_sc_hd__xnor2_1 _08062_ (.A(_01653_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__a21o_1 _08063_ (.A1(_01556_),
    .A2(_01659_),
    .B1(_01480_),
    .X(_01660_));
 sky130_fd_sc_hd__clkbuf_4 _08064_ (.A(_01512_),
    .X(_01661_));
 sky130_fd_sc_hd__o221a_1 _08065_ (.A1(_01539_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_01657_),
    .B2(_01660_),
    .C1(_01661_),
    .X(_00167_));
 sky130_fd_sc_hd__and2b_1 _08066_ (.A_N(net40),
    .B(net22),
    .X(_01662_));
 sky130_fd_sc_hd__and2b_1 _08067_ (.A_N(net22),
    .B(net40),
    .X(_01663_));
 sky130_fd_sc_hd__nor2_1 _08068_ (.A(_01662_),
    .B(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__and2_1 _08069_ (.A(net38),
    .B(net56),
    .X(_01665_));
 sky130_fd_sc_hd__o21ba_1 _08070_ (.A1(_01653_),
    .A2(_01655_),
    .B1_N(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__xnor2_1 _08071_ (.A(_01664_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__or2_1 _08072_ (.A(_01662_),
    .B(_01663_),
    .X(_01668_));
 sky130_fd_sc_hd__clkbuf_2 _08073_ (.A(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__or2b_1 _08074_ (.A(net56),
    .B_N(net38),
    .X(_01670_));
 sky130_fd_sc_hd__or2b_1 _08075_ (.A(net38),
    .B_N(net56),
    .X(_01671_));
 sky130_fd_sc_hd__nand2_2 _08076_ (.A(_01670_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__or2_1 _08077_ (.A(_01638_),
    .B(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__a21o_1 _08078_ (.A1(_01637_),
    .A2(_01671_),
    .B1(_01651_),
    .X(_01674_));
 sky130_fd_sc_hd__o21a_1 _08079_ (.A1(_01647_),
    .A2(_01673_),
    .B1(_01674_),
    .X(_01675_));
 sky130_fd_sc_hd__o21ai_1 _08080_ (.A1(_01669_),
    .A2(_01675_),
    .B1(_01470_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21o_1 _08081_ (.A1(_01669_),
    .A2(_01675_),
    .B1(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__o211ai_1 _08082_ (.A1(_01562_),
    .A2(_01667_),
    .B1(_01677_),
    .C1(_01485_),
    .Y(_01678_));
 sky130_fd_sc_hd__o211a_1 _08083_ (.A1(_01463_),
    .A2(net514),
    .B1(_01635_),
    .C1(_01678_),
    .X(_00168_));
 sky130_fd_sc_hd__and2b_1 _08084_ (.A_N(net41),
    .B(net23),
    .X(_01679_));
 sky130_fd_sc_hd__and2b_1 _08085_ (.A_N(net23),
    .B(net41),
    .X(_01680_));
 sky130_fd_sc_hd__nor2_2 _08086_ (.A(_01679_),
    .B(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(net22),
    .B(net40),
    .Y(_01682_));
 sky130_fd_sc_hd__o21a_1 _08088_ (.A1(_01664_),
    .A2(_01666_),
    .B1(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__xnor2_1 _08089_ (.A(_01681_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__nor2_1 _08090_ (.A(_01562_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__o21ba_1 _08091_ (.A1(_01669_),
    .A2(_01675_),
    .B1_N(_01663_),
    .X(_01686_));
 sky130_fd_sc_hd__xnor2_1 _08092_ (.A(_01681_),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__a21o_1 _08093_ (.A1(_01556_),
    .A2(_01687_),
    .B1(_01480_),
    .X(_01688_));
 sky130_fd_sc_hd__o221a_1 _08094_ (.A1(_01539_),
    .A2(net632),
    .B1(_01685_),
    .B2(_01688_),
    .C1(_01661_),
    .X(_00169_));
 sky130_fd_sc_hd__and2b_1 _08095_ (.A_N(net42),
    .B(net24),
    .X(_01689_));
 sky130_fd_sc_hd__and2b_1 _08096_ (.A_N(net24),
    .B(net42),
    .X(_01690_));
 sky130_fd_sc_hd__nor2_4 _08097_ (.A(_01689_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__o2111a_1 _08098_ (.A1(_01679_),
    .A2(_01680_),
    .B1(_01638_),
    .C1(_01672_),
    .D1(_01669_),
    .X(_01692_));
 sky130_fd_sc_hd__a21o_1 _08099_ (.A1(_01672_),
    .A2(_01654_),
    .B1(_01665_),
    .X(_01693_));
 sky130_fd_sc_hd__nand2_1 _08100_ (.A(_01669_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21oi_1 _08101_ (.A1(_01682_),
    .A2(_01694_),
    .B1(_01681_),
    .Y(_01695_));
 sky130_fd_sc_hd__a21o_1 _08102_ (.A1(net23),
    .A2(net41),
    .B1(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__a21oi_2 _08103_ (.A1(_01641_),
    .A2(_01692_),
    .B1(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__xnor2_1 _08104_ (.A(_01691_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__nor2_1 _08105_ (.A(_01562_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_2 _08106_ (.A(_01664_),
    .B(_01681_),
    .Y(_01700_));
 sky130_fd_sc_hd__inv_2 _08107_ (.A(_01679_),
    .Y(_01701_));
 sky130_fd_sc_hd__a21oi_1 _08108_ (.A1(_01663_),
    .A2(_01701_),
    .B1(_01680_),
    .Y(_01702_));
 sky130_fd_sc_hd__o21ai_2 _08109_ (.A1(_01675_),
    .A2(_01700_),
    .B1(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__xor2_1 _08110_ (.A(_01691_),
    .B(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__a21o_1 _08111_ (.A1(_01556_),
    .A2(_01704_),
    .B1(_01480_),
    .X(_01705_));
 sky130_fd_sc_hd__o221a_1 _08112_ (.A1(_01539_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_01699_),
    .B2(_01705_),
    .C1(_01661_),
    .X(_00170_));
 sky130_fd_sc_hd__nand2b_1 _08113_ (.A_N(net43),
    .B(net25),
    .Y(_01706_));
 sky130_fd_sc_hd__or2b_1 _08114_ (.A(net25),
    .B_N(net43),
    .X(_01707_));
 sky130_fd_sc_hd__nand2_1 _08115_ (.A(_01706_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__inv_2 _08116_ (.A(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _08117_ (.A(net24),
    .B(net42),
    .Y(_01710_));
 sky130_fd_sc_hd__o21a_1 _08118_ (.A1(_01691_),
    .A2(_01697_),
    .B1(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__xnor2_1 _08119_ (.A(_01709_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__nor2_1 _08120_ (.A(_01562_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__a21oi_1 _08121_ (.A1(_01691_),
    .A2(_01703_),
    .B1(_01690_),
    .Y(_01714_));
 sky130_fd_sc_hd__xnor2_1 _08122_ (.A(_01709_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__a21o_1 _08123_ (.A1(_01472_),
    .A2(_01715_),
    .B1(_01480_),
    .X(_01716_));
 sky130_fd_sc_hd__o221a_1 _08124_ (.A1(_01539_),
    .A2(net596),
    .B1(_01713_),
    .B2(_01716_),
    .C1(_01661_),
    .X(_00171_));
 sky130_fd_sc_hd__clkbuf_4 _08125_ (.A(_01457_),
    .X(_01717_));
 sky130_fd_sc_hd__inv_2 _08126_ (.A(net26),
    .Y(_01718_));
 sky130_fd_sc_hd__nor2_1 _08127_ (.A(_01718_),
    .B(net44),
    .Y(_01719_));
 sky130_fd_sc_hd__and2_1 _08128_ (.A(_01718_),
    .B(net44),
    .X(_01720_));
 sky130_fd_sc_hd__or2_1 _08129_ (.A(_01719_),
    .B(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__clkbuf_2 _08130_ (.A(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__nand2_1 _08131_ (.A(net25),
    .B(net43),
    .Y(_01723_));
 sky130_fd_sc_hd__o21ai_1 _08132_ (.A1(_01709_),
    .A2(_01710_),
    .B1(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__or3_1 _08133_ (.A(_01691_),
    .B(_01697_),
    .C(_01709_),
    .X(_01725_));
 sky130_fd_sc_hd__or2b_1 _08134_ (.A(_01724_),
    .B_N(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__xnor2_1 _08135_ (.A(_01722_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__and3_1 _08136_ (.A(_01691_),
    .B(_01706_),
    .C(_01707_),
    .X(_01728_));
 sky130_fd_sc_hd__and2b_1 _08137_ (.A_N(net25),
    .B(net43),
    .X(_01729_));
 sky130_fd_sc_hd__o21ai_1 _08138_ (.A1(_01690_),
    .A2(_01729_),
    .B1(_01706_),
    .Y(_01730_));
 sky130_fd_sc_hd__a21boi_1 _08139_ (.A1(_01703_),
    .A2(_01728_),
    .B1_N(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__nor2_1 _08140_ (.A(_01722_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__a21o_1 _08141_ (.A1(_01722_),
    .A2(_01731_),
    .B1(_01572_),
    .X(_01733_));
 sky130_fd_sc_hd__o221ai_1 _08142_ (.A1(_01556_),
    .A2(_01727_),
    .B1(_01732_),
    .B2(_01733_),
    .C1(_01485_),
    .Y(_01734_));
 sky130_fd_sc_hd__o211a_1 _08143_ (.A1(_01717_),
    .A2(net410),
    .B1(_01635_),
    .C1(_01734_),
    .X(_00172_));
 sky130_fd_sc_hd__and2b_1 _08144_ (.A_N(net27),
    .B(net45),
    .X(_01735_));
 sky130_fd_sc_hd__or2b_1 _08145_ (.A(net45),
    .B_N(net27),
    .X(_01736_));
 sky130_fd_sc_hd__and2b_1 _08146_ (.A_N(_01735_),
    .B(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__buf_2 _08147_ (.A(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__o21ba_1 _08148_ (.A1(_01722_),
    .A2(_01731_),
    .B1_N(_01720_),
    .X(_01739_));
 sky130_fd_sc_hd__xnor2_1 _08149_ (.A(_01738_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _08150_ (.A(net26),
    .B(net44),
    .Y(_01741_));
 sky130_fd_sc_hd__a21bo_1 _08151_ (.A1(_01722_),
    .A2(_01726_),
    .B1_N(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__xor2_1 _08152_ (.A(_01738_),
    .B(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__nor2_1 _08153_ (.A(_01472_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__a211o_1 _08154_ (.A1(_01556_),
    .A2(_01740_),
    .B1(_01744_),
    .C1(_01454_),
    .X(_01745_));
 sky130_fd_sc_hd__o211a_1 _08155_ (.A1(_01717_),
    .A2(net446),
    .B1(_01635_),
    .C1(_01745_),
    .X(_00173_));
 sky130_fd_sc_hd__and2b_1 _08156_ (.A_N(net46),
    .B(net28),
    .X(_01746_));
 sky130_fd_sc_hd__and2b_1 _08157_ (.A_N(net28),
    .B(net46),
    .X(_01747_));
 sky130_fd_sc_hd__or2_2 _08158_ (.A(_01746_),
    .B(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__inv_2 _08159_ (.A(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_2 _08160_ (.A(_01719_),
    .B(_01720_),
    .Y(_01750_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(_01722_),
    .B(_01724_),
    .Y(_01751_));
 sky130_fd_sc_hd__a21oi_1 _08162_ (.A1(_01741_),
    .A2(_01751_),
    .B1(_01738_),
    .Y(_01752_));
 sky130_fd_sc_hd__a21oi_1 _08163_ (.A1(net27),
    .A2(net45),
    .B1(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__o31a_1 _08164_ (.A1(_01750_),
    .A2(_01725_),
    .A3(_01738_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__xnor2_1 _08165_ (.A(_01749_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__and2_1 _08166_ (.A(_01750_),
    .B(_01738_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(_01728_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__inv_2 _08168_ (.A(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__nand2_1 _08169_ (.A(_01750_),
    .B(_01738_),
    .Y(_01759_));
 sky130_fd_sc_hd__o2bb2a_1 _08170_ (.A1_N(_01703_),
    .A2_N(_01758_),
    .B1(_01759_),
    .B2(_01730_),
    .X(_01760_));
 sky130_fd_sc_hd__a21oi_1 _08171_ (.A1(_01720_),
    .A2(_01736_),
    .B1(_01735_),
    .Y(_01761_));
 sky130_fd_sc_hd__a21oi_1 _08172_ (.A1(_01760_),
    .A2(_01761_),
    .B1(_01748_),
    .Y(_01762_));
 sky130_fd_sc_hd__a31o_1 _08173_ (.A1(_01748_),
    .A2(_01760_),
    .A3(_01761_),
    .B1(_01329_),
    .X(_01763_));
 sky130_fd_sc_hd__o221a_1 _08174_ (.A1(_01472_),
    .A2(_01755_),
    .B1(_01762_),
    .B2(_01763_),
    .C1(_01457_),
    .X(_01764_));
 sky130_fd_sc_hd__buf_4 _08175_ (.A(_01251_),
    .X(_01765_));
 sky130_fd_sc_hd__clkbuf_8 _08176_ (.A(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__o21ai_1 _08177_ (.A1(_01529_),
    .A2(net454),
    .B1(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _08178_ (.A(_01764_),
    .B(_01767_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _08179_ (.A(net28),
    .B(net46),
    .Y(_01768_));
 sky130_fd_sc_hd__o21ai_1 _08180_ (.A1(_01749_),
    .A2(_01754_),
    .B1(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__xor2_2 _08181_ (.A(net29),
    .B(net47),
    .X(_01770_));
 sky130_fd_sc_hd__xnor2_1 _08182_ (.A(_01769_),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _08183_ (.A(_01556_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__or3_1 _08184_ (.A(_01747_),
    .B(_01762_),
    .C(_01770_),
    .X(_01773_));
 sky130_fd_sc_hd__o21ai_1 _08185_ (.A1(_01747_),
    .A2(_01762_),
    .B1(_01770_),
    .Y(_01774_));
 sky130_fd_sc_hd__a21oi_1 _08186_ (.A1(_01773_),
    .A2(_01774_),
    .B1(_01330_),
    .Y(_01775_));
 sky130_fd_sc_hd__or2_1 _08187_ (.A(_01464_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[17] ),
    .X(_01776_));
 sky130_fd_sc_hd__o311a_1 _08188_ (.A1(_01454_),
    .A2(_01772_),
    .A3(_01775_),
    .B1(_01776_),
    .C1(_01766_),
    .X(_00175_));
 sky130_fd_sc_hd__and2_1 _08189_ (.A(net39),
    .B(_01329_),
    .X(_01777_));
 sky130_fd_sc_hd__nor2_1 _08190_ (.A(_01559_),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__a21o_1 _08191_ (.A1(_01559_),
    .A2(_01777_),
    .B1(_01453_),
    .X(_01779_));
 sky130_fd_sc_hd__o221a_1 _08192_ (.A1(_01539_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .B1(_01778_),
    .B2(_01779_),
    .C1(_01661_),
    .X(_00176_));
 sky130_fd_sc_hd__o21ai_1 _08193_ (.A1(_01553_),
    .A2(_01570_),
    .B1(_01569_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _08194_ (.A(_01565_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__and2_1 _08195_ (.A(_01565_),
    .B(_01780_),
    .X(_01782_));
 sky130_fd_sc_hd__o31a_1 _08196_ (.A1(_01470_),
    .A2(_01781_),
    .A3(_01782_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ),
    .X(_01783_));
 sky130_fd_sc_hd__o21ai_2 _08197_ (.A1(_01330_),
    .A2(_01568_),
    .B1(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o211a_1 _08198_ (.A1(_01717_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_01635_),
    .C1(_01784_),
    .X(_00177_));
 sky130_fd_sc_hd__nor2_1 _08199_ (.A(_01563_),
    .B(_01782_),
    .Y(_01785_));
 sky130_fd_sc_hd__xnor2_1 _08200_ (.A(_01579_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__mux2_1 _08201_ (.A0(_01582_),
    .A1(_01786_),
    .S(_01329_),
    .X(_01787_));
 sky130_fd_sc_hd__nand2_1 _08202_ (.A(_01465_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__o211a_1 _08203_ (.A1(_01717_),
    .A2(net631),
    .B1(_01635_),
    .C1(_01788_),
    .X(_00178_));
 sky130_fd_sc_hd__nand2_1 _08204_ (.A(_01565_),
    .B(_01780_),
    .Y(_01789_));
 sky130_fd_sc_hd__a31o_1 _08205_ (.A1(_01577_),
    .A2(_01584_),
    .A3(_01789_),
    .B1(_01576_),
    .X(_01790_));
 sky130_fd_sc_hd__nor2_1 _08206_ (.A(_01589_),
    .B(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__a21o_1 _08207_ (.A1(_01589_),
    .A2(_01790_),
    .B1(_01470_),
    .X(_01792_));
 sky130_fd_sc_hd__o221a_1 _08208_ (.A1(_01572_),
    .A2(_01592_),
    .B1(_01791_),
    .B2(_01792_),
    .C1(_01457_),
    .X(_01793_));
 sky130_fd_sc_hd__buf_6 _08209_ (.A(_01765_),
    .X(_01794_));
 sky130_fd_sc_hd__o21ai_1 _08210_ (.A1(_01529_),
    .A2(net542),
    .B1(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _08211_ (.A(_01793_),
    .B(_01795_),
    .Y(_00179_));
 sky130_fd_sc_hd__o21ai_1 _08212_ (.A1(_01589_),
    .A2(_01790_),
    .B1(_01587_),
    .Y(_01796_));
 sky130_fd_sc_hd__xnor2_1 _08213_ (.A(_01599_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__mux2_1 _08214_ (.A0(_01602_),
    .A1(_01797_),
    .S(_01329_),
    .X(_01798_));
 sky130_fd_sc_hd__nand2_1 _08215_ (.A(_01465_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__o211a_1 _08216_ (.A1(_01717_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .B1(_01635_),
    .C1(_01799_),
    .X(_00180_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_01597_),
    .B(_01796_),
    .Y(_01800_));
 sky130_fd_sc_hd__a21oi_1 _08218_ (.A1(_01598_),
    .A2(_01800_),
    .B1(_01612_),
    .Y(_01801_));
 sky130_fd_sc_hd__a31o_1 _08219_ (.A1(_01598_),
    .A2(_01612_),
    .A3(_01800_),
    .B1(_01470_),
    .X(_01802_));
 sky130_fd_sc_hd__o221a_1 _08220_ (.A1(_01572_),
    .A2(_01621_),
    .B1(_01801_),
    .B2(_01802_),
    .C1(_01457_),
    .X(_01803_));
 sky130_fd_sc_hd__o21ai_1 _08221_ (.A1(_01529_),
    .A2(net508),
    .B1(_01794_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _08222_ (.A(_01803_),
    .B(_01804_),
    .Y(_00181_));
 sky130_fd_sc_hd__o21ai_1 _08223_ (.A1(_01609_),
    .A2(_01801_),
    .B1(_01627_),
    .Y(_01805_));
 sky130_fd_sc_hd__or3_1 _08224_ (.A(_01609_),
    .B(_01627_),
    .C(_01801_),
    .X(_01806_));
 sky130_fd_sc_hd__a21oi_1 _08225_ (.A1(_01805_),
    .A2(_01806_),
    .B1(_01562_),
    .Y(_01807_));
 sky130_fd_sc_hd__o21ai_1 _08226_ (.A1(_01330_),
    .A2(_01630_),
    .B1(_01529_),
    .Y(_01808_));
 sky130_fd_sc_hd__o221a_1 _08227_ (.A1(_01465_),
    .A2(net511),
    .B1(_01807_),
    .B2(_01808_),
    .C1(_01661_),
    .X(_00182_));
 sky130_fd_sc_hd__and3_1 _08228_ (.A(_01599_),
    .B(_01643_),
    .C(_01791_),
    .X(_01809_));
 sky130_fd_sc_hd__a21oi_2 _08229_ (.A1(_01625_),
    .A2(_01646_),
    .B1(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_01638_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__a21o_1 _08231_ (.A1(_01638_),
    .A2(_01810_),
    .B1(_01472_),
    .X(_01812_));
 sky130_fd_sc_hd__o221ai_4 _08232_ (.A1(_01330_),
    .A2(_01642_),
    .B1(_01811_),
    .B2(_01812_),
    .C1(_01485_),
    .Y(_01813_));
 sky130_fd_sc_hd__o211a_1 _08233_ (.A1(_01717_),
    .A2(net309),
    .B1(_01635_),
    .C1(_01813_),
    .X(_00183_));
 sky130_fd_sc_hd__o21a_1 _08234_ (.A1(_01638_),
    .A2(_01810_),
    .B1(_01636_),
    .X(_01814_));
 sky130_fd_sc_hd__xnor2_1 _08235_ (.A(_01672_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__mux2_1 _08236_ (.A0(_01656_),
    .A1(_01815_),
    .S(_01329_),
    .X(_01816_));
 sky130_fd_sc_hd__nand2_1 _08237_ (.A(_01465_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__o211a_1 _08238_ (.A1(_01717_),
    .A2(net458),
    .B1(_01635_),
    .C1(_01817_),
    .X(_00184_));
 sky130_fd_sc_hd__a21o_1 _08239_ (.A1(_01636_),
    .A2(_01670_),
    .B1(_01652_),
    .X(_01818_));
 sky130_fd_sc_hd__o21a_1 _08240_ (.A1(_01673_),
    .A2(_01810_),
    .B1(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__nor2_1 _08241_ (.A(_01669_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__a21o_1 _08242_ (.A1(_01669_),
    .A2(_01819_),
    .B1(_01472_),
    .X(_01821_));
 sky130_fd_sc_hd__o221ai_2 _08243_ (.A1(_01572_),
    .A2(_01667_),
    .B1(_01820_),
    .B2(_01821_),
    .C1(_01485_),
    .Y(_01822_));
 sky130_fd_sc_hd__o211a_1 _08244_ (.A1(_01717_),
    .A2(net475),
    .B1(_01635_),
    .C1(_01822_),
    .X(_00185_));
 sky130_fd_sc_hd__clkbuf_4 _08245_ (.A(_01455_),
    .X(_01823_));
 sky130_fd_sc_hd__or2_1 _08246_ (.A(_01662_),
    .B(_01820_),
    .X(_01824_));
 sky130_fd_sc_hd__xnor2_1 _08247_ (.A(_01681_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__mux2_1 _08248_ (.A0(_01684_),
    .A1(_01825_),
    .S(_01329_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _08249_ (.A(_01465_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__o211a_1 _08250_ (.A1(_01717_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_01823_),
    .C1(_01827_),
    .X(_00186_));
 sky130_fd_sc_hd__nor2_1 _08251_ (.A(_01330_),
    .B(_01698_),
    .Y(_01828_));
 sky130_fd_sc_hd__or2b_1 _08252_ (.A(_01680_),
    .B_N(_01662_),
    .X(_01829_));
 sky130_fd_sc_hd__o211ai_4 _08253_ (.A1(_01700_),
    .A2(_01819_),
    .B1(_01829_),
    .C1(_01701_),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _08254_ (.A(_01691_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__a21o_1 _08255_ (.A1(_01691_),
    .A2(_01830_),
    .B1(_01470_),
    .X(_01832_));
 sky130_fd_sc_hd__o21ai_1 _08256_ (.A1(_01831_),
    .A2(_01832_),
    .B1(_01529_),
    .Y(_01833_));
 sky130_fd_sc_hd__o221a_1 _08257_ (.A1(_01465_),
    .A2(net630),
    .B1(_01828_),
    .B2(_01833_),
    .C1(_01661_),
    .X(_00187_));
 sky130_fd_sc_hd__a21o_1 _08258_ (.A1(_01691_),
    .A2(_01830_),
    .B1(_01689_),
    .X(_01834_));
 sky130_fd_sc_hd__xnor2_1 _08259_ (.A(_01709_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_1 _08260_ (.A(_01562_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__o21ai_1 _08261_ (.A1(_01330_),
    .A2(_01712_),
    .B1(_01529_),
    .Y(_01837_));
 sky130_fd_sc_hd__o221a_1 _08262_ (.A1(_01465_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_01836_),
    .B2(_01837_),
    .C1(_01661_),
    .X(_00188_));
 sky130_fd_sc_hd__or2b_1 _08263_ (.A(net42),
    .B_N(net24),
    .X(_01838_));
 sky130_fd_sc_hd__a21oi_1 _08264_ (.A1(_01838_),
    .A2(_01706_),
    .B1(_01729_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21o_1 _08265_ (.A1(_01728_),
    .A2(_01830_),
    .B1(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__nor2_1 _08266_ (.A(_01750_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__a21o_1 _08267_ (.A1(_01750_),
    .A2(_01840_),
    .B1(_01470_),
    .X(_01842_));
 sky130_fd_sc_hd__o221a_1 _08268_ (.A1(_01572_),
    .A2(_01727_),
    .B1(_01841_),
    .B2(_01842_),
    .C1(_01457_),
    .X(_01843_));
 sky130_fd_sc_hd__o21ai_1 _08269_ (.A1(_01529_),
    .A2(net551),
    .B1(_01794_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _08270_ (.A(_01843_),
    .B(_01844_),
    .Y(_00189_));
 sky130_fd_sc_hd__a21oi_1 _08271_ (.A1(_01750_),
    .A2(_01840_),
    .B1(_01719_),
    .Y(_01845_));
 sky130_fd_sc_hd__xnor2_1 _08272_ (.A(_01738_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _08273_ (.A(_01572_),
    .B(_01743_),
    .Y(_01847_));
 sky130_fd_sc_hd__a211o_1 _08274_ (.A1(_01572_),
    .A2(_01846_),
    .B1(_01847_),
    .C1(_01454_),
    .X(_01848_));
 sky130_fd_sc_hd__o211a_1 _08275_ (.A1(_01717_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_01823_),
    .C1(_01848_),
    .X(_00190_));
 sky130_fd_sc_hd__nor2_1 _08276_ (.A(_01330_),
    .B(_01755_),
    .Y(_01849_));
 sky130_fd_sc_hd__a22oi_2 _08277_ (.A1(_01758_),
    .A2(_01830_),
    .B1(_01839_),
    .B2(_01756_),
    .Y(_01850_));
 sky130_fd_sc_hd__o31a_1 _08278_ (.A1(_01718_),
    .A2(net44),
    .A3(_01735_),
    .B1(_01736_),
    .X(_01851_));
 sky130_fd_sc_hd__a21oi_1 _08279_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_01748_),
    .Y(_01852_));
 sky130_fd_sc_hd__a31o_1 _08280_ (.A1(_01748_),
    .A2(_01850_),
    .A3(_01851_),
    .B1(_01472_),
    .X(_01853_));
 sky130_fd_sc_hd__nor2_1 _08281_ (.A(_01852_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__or2_1 _08282_ (.A(_01464_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ),
    .X(_01855_));
 sky130_fd_sc_hd__o311a_1 _08283_ (.A1(_01454_),
    .A2(_01849_),
    .A3(_01854_),
    .B1(_01855_),
    .C1(_01766_),
    .X(_00191_));
 sky130_fd_sc_hd__nor2_1 _08284_ (.A(_01330_),
    .B(_01771_),
    .Y(_01856_));
 sky130_fd_sc_hd__or3_1 _08285_ (.A(_01746_),
    .B(_01770_),
    .C(_01852_),
    .X(_01857_));
 sky130_fd_sc_hd__o21ai_1 _08286_ (.A1(_01746_),
    .A2(_01852_),
    .B1(_01770_),
    .Y(_01858_));
 sky130_fd_sc_hd__a21oi_1 _08287_ (.A1(_01857_),
    .A2(_01858_),
    .B1(_01562_),
    .Y(_01859_));
 sky130_fd_sc_hd__or2_1 _08288_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[17] ),
    .B(_01464_),
    .X(_01860_));
 sky130_fd_sc_hd__o311a_1 _08289_ (.A1(_01454_),
    .A2(_01856_),
    .A3(_01859_),
    .B1(_01860_),
    .C1(_01766_),
    .X(_00192_));
 sky130_fd_sc_hd__clkbuf_4 _08290_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_01861_));
 sky130_fd_sc_hd__clkbuf_4 _08291_ (.A(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__and2_1 _08292_ (.A(_01862_),
    .B(_01253_),
    .X(_01863_));
 sky130_fd_sc_hd__clkbuf_1 _08293_ (.A(_01863_),
    .X(_00193_));
 sky130_fd_sc_hd__inv_2 _08294_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_out ),
    .Y(_01864_));
 sky130_fd_sc_hd__clkbuf_4 _08295_ (.A(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__clkbuf_4 _08296_ (.A(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__buf_4 _08297_ (.A(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__clkbuf_4 _08298_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_out ),
    .X(_01868_));
 sky130_fd_sc_hd__clkbuf_4 _08299_ (.A(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__clkbuf_4 _08300_ (.A(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__or2_1 _08301_ (.A(net155),
    .B(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__o211a_1 _08302_ (.A1(_01867_),
    .A2(net203),
    .B1(_01823_),
    .C1(_01871_),
    .X(_00194_));
 sky130_fd_sc_hd__or2_1 _08303_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_01870_),
    .X(_01872_));
 sky130_fd_sc_hd__o211a_1 _08304_ (.A1(_01867_),
    .A2(net159),
    .B1(_01823_),
    .C1(_01872_),
    .X(_00195_));
 sky130_fd_sc_hd__buf_2 _08305_ (.A(_01868_),
    .X(_01873_));
 sky130_fd_sc_hd__or2_1 _08306_ (.A(net147),
    .B(_01873_),
    .X(_01874_));
 sky130_fd_sc_hd__o211a_1 _08307_ (.A1(_01867_),
    .A2(net165),
    .B1(_01823_),
    .C1(_01874_),
    .X(_00196_));
 sky130_fd_sc_hd__or2_1 _08308_ (.A(_01870_),
    .B(net650),
    .X(_01875_));
 sky130_fd_sc_hd__o211a_1 _08309_ (.A1(_01867_),
    .A2(net164),
    .B1(_01823_),
    .C1(_01875_),
    .X(_00197_));
 sky130_fd_sc_hd__clkbuf_4 _08310_ (.A(_01869_),
    .X(_01876_));
 sky130_fd_sc_hd__clkbuf_4 _08311_ (.A(_01869_),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_1 _08312_ (.A(_01877_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .Y(_01878_));
 sky130_fd_sc_hd__o211a_1 _08313_ (.A1(_01876_),
    .A2(net307),
    .B1(_01823_),
    .C1(_01878_),
    .X(_00198_));
 sky130_fd_sc_hd__inv_2 _08314_ (.A(_01549_),
    .Y(_01879_));
 sky130_fd_sc_hd__clkbuf_4 _08315_ (.A(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__buf_2 _08316_ (.A(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__buf_4 _08317_ (.A(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__xor2_2 _08318_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(_01883_));
 sky130_fd_sc_hd__xnor2_1 _08319_ (.A(_01882_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__or2_1 _08320_ (.A(_01873_),
    .B(net618),
    .X(_01885_));
 sky130_fd_sc_hd__o211a_1 _08321_ (.A1(_01867_),
    .A2(_01884_),
    .B1(_01885_),
    .C1(_01552_),
    .X(_00199_));
 sky130_fd_sc_hd__o21ai_1 _08322_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ),
    .Y(_01886_));
 sky130_fd_sc_hd__or3_1 _08323_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ),
    .C(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(_01887_));
 sky130_fd_sc_hd__o211a_1 _08324_ (.A1(_01550_),
    .A2(_01883_),
    .B1(_01886_),
    .C1(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__a211o_1 _08325_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01550_),
    .C1(_01883_),
    .X(_01889_));
 sky130_fd_sc_hd__nand2_1 _08326_ (.A(_01877_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__o221a_1 _08327_ (.A1(_01876_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B1(_01888_),
    .B2(_01890_),
    .C1(_01661_),
    .X(_00200_));
 sky130_fd_sc_hd__clkbuf_4 _08328_ (.A(_01869_),
    .X(_01891_));
 sky130_fd_sc_hd__o21a_1 _08329_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(_01892_));
 sky130_fd_sc_hd__a21oi_1 _08330_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ),
    .Y(_01893_));
 sky130_fd_sc_hd__mux2_1 _08331_ (.A0(_01892_),
    .A1(_01893_),
    .S(_01882_),
    .X(_01894_));
 sky130_fd_sc_hd__and2_1 _08332_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__o21ai_1 _08333_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(_01894_),
    .B1(_01877_),
    .Y(_01896_));
 sky130_fd_sc_hd__o221a_1 _08334_ (.A1(_01891_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B1(_01895_),
    .B2(_01896_),
    .C1(_01661_),
    .X(_00201_));
 sky130_fd_sc_hd__or2_1 _08335_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_01892_),
    .X(_01897_));
 sky130_fd_sc_hd__and2b_1 _08336_ (.A_N(_01893_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(_01898_));
 sky130_fd_sc_hd__nor2_1 _08337_ (.A(_01550_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__a21oi_1 _08338_ (.A1(_01550_),
    .A2(_01897_),
    .B1(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__o21ai_1 _08339_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_01900_),
    .B1(_01869_),
    .Y(_01901_));
 sky130_fd_sc_hd__a21o_1 _08340_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_01900_),
    .B1(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__o211a_1 _08341_ (.A1(_01876_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B1(_01823_),
    .C1(_01902_),
    .X(_00202_));
 sky130_fd_sc_hd__o21a_1 _08342_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_01898_),
    .B1(_01882_),
    .X(_01903_));
 sky130_fd_sc_hd__a21oi_1 _08343_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_01897_),
    .B1(_01882_),
    .Y(_01904_));
 sky130_fd_sc_hd__inv_2 _08344_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_01905_));
 sky130_fd_sc_hd__o21a_1 _08345_ (.A1(_01903_),
    .A2(_01904_),
    .B1(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__o31ai_1 _08346_ (.A1(_01905_),
    .A2(_01903_),
    .A3(_01904_),
    .B1(_01870_),
    .Y(_01907_));
 sky130_fd_sc_hd__clkbuf_4 _08347_ (.A(_01512_),
    .X(_01908_));
 sky130_fd_sc_hd__o221a_1 _08348_ (.A1(_01891_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B1(_01906_),
    .B2(_01907_),
    .C1(_01908_),
    .X(_00203_));
 sky130_fd_sc_hd__inv_2 _08349_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[8] ),
    .Y(_01909_));
 sky130_fd_sc_hd__a21oi_1 _08350_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_01897_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_01910_));
 sky130_fd_sc_hd__a22o_1 _08351_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(_01903_),
    .B1(_01910_),
    .B2(_01550_),
    .X(_01911_));
 sky130_fd_sc_hd__a21oi_1 _08352_ (.A1(_01909_),
    .A2(_01911_),
    .B1(_01866_),
    .Y(_01912_));
 sky130_fd_sc_hd__o21ai_1 _08353_ (.A1(_01909_),
    .A2(_01911_),
    .B1(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__o211a_1 _08354_ (.A1(_01876_),
    .A2(net398),
    .B1(_01823_),
    .C1(_01913_),
    .X(_00204_));
 sky130_fd_sc_hd__o211a_1 _08355_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_01898_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[8] ),
    .C1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(_01914_));
 sky130_fd_sc_hd__nor2_1 _08356_ (.A(_01550_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _08357_ (.A(_01909_),
    .B(_01910_),
    .Y(_01916_));
 sky130_fd_sc_hd__and2_1 _08358_ (.A(_01550_),
    .B(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__inv_2 _08359_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_01918_));
 sky130_fd_sc_hd__o21a_1 _08360_ (.A1(_01915_),
    .A2(_01917_),
    .B1(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__o31ai_1 _08361_ (.A1(_01918_),
    .A2(_01915_),
    .A3(_01917_),
    .B1(_01870_),
    .Y(_01920_));
 sky130_fd_sc_hd__o221a_1 _08362_ (.A1(_01891_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_01919_),
    .B2(_01920_),
    .C1(_01908_),
    .X(_00205_));
 sky130_fd_sc_hd__a2bb2o_1 _08363_ (.A1_N(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2_N(_01914_),
    .B1(_01916_),
    .B2(_01550_),
    .X(_01921_));
 sky130_fd_sc_hd__nand2_1 _08364_ (.A(_01550_),
    .B(_01918_),
    .Y(_01922_));
 sky130_fd_sc_hd__a21oi_1 _08365_ (.A1(_01921_),
    .A2(_01922_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ),
    .Y(_01923_));
 sky130_fd_sc_hd__clkbuf_4 _08366_ (.A(_01865_),
    .X(_01924_));
 sky130_fd_sc_hd__a31o_1 _08367_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_01921_),
    .A3(_01922_),
    .B1(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__o221a_1 _08368_ (.A1(_01891_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_01923_),
    .B2(_01925_),
    .C1(_01908_),
    .X(_00206_));
 sky130_fd_sc_hd__inv_2 _08369_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[11] ),
    .Y(_01926_));
 sky130_fd_sc_hd__a21oi_1 _08370_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_01916_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ),
    .Y(_01927_));
 sky130_fd_sc_hd__o21a_1 _08371_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_01914_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _08372_ (.A0(_01927_),
    .A1(_01928_),
    .S(_01882_),
    .X(_01929_));
 sky130_fd_sc_hd__and2_1 _08373_ (.A(_01926_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__o21ai_1 _08374_ (.A1(_01926_),
    .A2(_01929_),
    .B1(_01877_),
    .Y(_01931_));
 sky130_fd_sc_hd__o221a_1 _08375_ (.A1(_01891_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B1(_01930_),
    .B2(_01931_),
    .C1(_01908_),
    .X(_00207_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(_01926_),
    .B(_01927_),
    .Y(_01932_));
 sky130_fd_sc_hd__and2_1 _08377_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_01928_),
    .X(_01933_));
 sky130_fd_sc_hd__inv_2 _08378_ (.A(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__mux2_1 _08379_ (.A0(_01932_),
    .A1(_01934_),
    .S(_01882_),
    .X(_01935_));
 sky130_fd_sc_hd__and2_1 _08380_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__o21ai_1 _08381_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_01935_),
    .B1(_01870_),
    .Y(_01937_));
 sky130_fd_sc_hd__o221a_1 _08382_ (.A1(_01891_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_01936_),
    .B2(_01937_),
    .C1(_01908_),
    .X(_00208_));
 sky130_fd_sc_hd__a31o_1 _08383_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(_01928_),
    .B1(_01549_),
    .X(_01938_));
 sky130_fd_sc_hd__o21ai_1 _08384_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_01932_),
    .B1(_01549_),
    .Y(_01939_));
 sky130_fd_sc_hd__a21oi_1 _08385_ (.A1(_01938_),
    .A2(_01939_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ),
    .Y(_01940_));
 sky130_fd_sc_hd__a31o_1 _08386_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_01938_),
    .A3(_01939_),
    .B1(_01924_),
    .X(_01941_));
 sky130_fd_sc_hd__o221a_1 _08387_ (.A1(_01891_),
    .A2(net628),
    .B1(_01940_),
    .B2(_01941_),
    .C1(_01908_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _08388_ (.A0(_01938_),
    .A1(_01939_),
    .S(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(_01942_));
 sky130_fd_sc_hd__a21oi_1 _08389_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_01942_),
    .B1(_01866_),
    .Y(_01943_));
 sky130_fd_sc_hd__o21ai_1 _08390_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_01942_),
    .B1(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__o211a_1 _08391_ (.A1(_01876_),
    .A2(net481),
    .B1(_01823_),
    .C1(_01944_),
    .X(_00210_));
 sky130_fd_sc_hd__clkbuf_4 _08392_ (.A(_01455_),
    .X(_01945_));
 sky130_fd_sc_hd__o211a_1 _08393_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_01932_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ),
    .C1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(_01946_));
 sky130_fd_sc_hd__a211o_1 _08394_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_01933_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ),
    .C1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(_01947_));
 sky130_fd_sc_hd__inv_2 _08395_ (.A(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__mux2_1 _08396_ (.A0(_01946_),
    .A1(_01948_),
    .S(_01882_),
    .X(_01949_));
 sky130_fd_sc_hd__xnor2_1 _08397_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__nand2_1 _08398_ (.A(_01877_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__o211a_1 _08399_ (.A1(_01876_),
    .A2(net427),
    .B1(_01945_),
    .C1(_01951_),
    .X(_00211_));
 sky130_fd_sc_hd__o21a_1 _08400_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_01947_),
    .B1(_01882_),
    .X(_01952_));
 sky130_fd_sc_hd__a21oi_1 _08401_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_01946_),
    .B1(_01882_),
    .Y(_01953_));
 sky130_fd_sc_hd__o21a_1 _08402_ (.A1(_01952_),
    .A2(_01953_),
    .B1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_01954_));
 sky130_fd_sc_hd__o31ai_1 _08403_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_01952_),
    .A3(_01953_),
    .B1(_01870_),
    .Y(_01955_));
 sky130_fd_sc_hd__o221a_1 _08404_ (.A1(_01891_),
    .A2(net531),
    .B1(_01954_),
    .B2(_01955_),
    .C1(_01908_),
    .X(_00212_));
 sky130_fd_sc_hd__inv_2 _08405_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[16] ),
    .Y(_01956_));
 sky130_fd_sc_hd__o21ba_1 _08406_ (.A1(_01956_),
    .A2(_01953_),
    .B1_N(_01952_),
    .X(_01957_));
 sky130_fd_sc_hd__clkbuf_4 _08407_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_01958_));
 sky130_fd_sc_hd__buf_2 _08408_ (.A(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__or2_1 _08409_ (.A(_01873_),
    .B(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__o211a_1 _08410_ (.A1(_01867_),
    .A2(_01957_),
    .B1(_01960_),
    .C1(_01552_),
    .X(_00213_));
 sky130_fd_sc_hd__inv_2 _08411_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .Y(_01961_));
 sky130_fd_sc_hd__nor2_1 _08412_ (.A(_01961_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ),
    .Y(_01962_));
 sky130_fd_sc_hd__a21o_1 _08413_ (.A1(_01961_),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ),
    .B1(_01866_),
    .X(_01963_));
 sky130_fd_sc_hd__o221a_1 _08414_ (.A1(_01891_),
    .A2(net465),
    .B1(_01962_),
    .B2(_01963_),
    .C1(_01908_),
    .X(_00214_));
 sky130_fd_sc_hd__and2b_1 _08415_ (.A_N(_01549_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .X(_01964_));
 sky130_fd_sc_hd__xnor2_1 _08416_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__xnor2_1 _08417_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__xor2_1 _08418_ (.A(_01962_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__or2_1 _08419_ (.A(_01873_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_01968_));
 sky130_fd_sc_hd__o211a_1 _08420_ (.A1(_01867_),
    .A2(_01967_),
    .B1(_01968_),
    .C1(_01552_),
    .X(_00215_));
 sky130_fd_sc_hd__and2_1 _08421_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B(_01965_),
    .X(_01969_));
 sky130_fd_sc_hd__nor2_1 _08422_ (.A(_01962_),
    .B(_01966_),
    .Y(_01970_));
 sky130_fd_sc_hd__o21ba_1 _08423_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .B1_N(_01549_),
    .X(_01971_));
 sky130_fd_sc_hd__xnor2_1 _08424_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__or2_1 _08425_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__nand2_1 _08426_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .B(_01972_),
    .Y(_01974_));
 sky130_fd_sc_hd__and2_1 _08427_ (.A(_01973_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__o21ai_2 _08428_ (.A1(_01969_),
    .A2(_01970_),
    .B1(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__o31a_1 _08429_ (.A1(_01969_),
    .A2(_01970_),
    .A3(_01975_),
    .B1(_01868_),
    .X(_01977_));
 sky130_fd_sc_hd__a22oi_1 _08430_ (.A1(_01865_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_01976_),
    .B2(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__buf_4 _08431_ (.A(_01251_),
    .X(_01979_));
 sky130_fd_sc_hd__and2b_1 _08432_ (.A_N(_01978_),
    .B(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__clkbuf_1 _08433_ (.A(_01980_),
    .X(_00216_));
 sky130_fd_sc_hd__clkbuf_4 _08434_ (.A(_01765_),
    .X(_01981_));
 sky130_fd_sc_hd__o31a_1 _08435_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ),
    .A3(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .B1(_01879_),
    .X(_01982_));
 sky130_fd_sc_hd__xnor2_1 _08436_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[4] ),
    .B(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _08437_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__or2_1 _08438_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ),
    .B(_01983_),
    .X(_01985_));
 sky130_fd_sc_hd__and2_1 _08439_ (.A(_01984_),
    .B(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__nand2_1 _08440_ (.A(_01974_),
    .B(_01976_),
    .Y(_01987_));
 sky130_fd_sc_hd__xor2_1 _08441_ (.A(_01986_),
    .B(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _08442_ (.A0(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_01988_),
    .S(_01868_),
    .X(_01989_));
 sky130_fd_sc_hd__and2_1 _08443_ (.A(_01981_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__clkbuf_1 _08444_ (.A(_01990_),
    .X(_00217_));
 sky130_fd_sc_hd__a21bo_1 _08445_ (.A1(_01974_),
    .A2(_01976_),
    .B1_N(_01986_),
    .X(_01991_));
 sky130_fd_sc_hd__or4_2 _08446_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[4] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ),
    .C(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ),
    .D(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .X(_01992_));
 sky130_fd_sc_hd__nand2_1 _08447_ (.A(_01880_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__xor2_1 _08448_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .B(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__or2_1 _08450_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ),
    .B(_01994_),
    .X(_01996_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_01995_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__a21oi_4 _08452_ (.A1(_01984_),
    .A2(_01991_),
    .B1(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__and3_1 _08453_ (.A(_01984_),
    .B(_01991_),
    .C(_01997_),
    .X(_01999_));
 sky130_fd_sc_hd__o21ai_1 _08454_ (.A1(_01998_),
    .A2(_01999_),
    .B1(_01877_),
    .Y(_02000_));
 sky130_fd_sc_hd__o211a_1 _08455_ (.A1(_01876_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B1(_01945_),
    .C1(_02000_),
    .X(_00218_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_01998_),
    .Y(_02001_));
 sky130_fd_sc_hd__inv_2 _08457_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_02002_));
 sky130_fd_sc_hd__o21a_1 _08458_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .A2(_01992_),
    .B1(_01880_),
    .X(_02003_));
 sky130_fd_sc_hd__xnor2_4 _08459_ (.A(_02002_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__xnor2_4 _08460_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ),
    .B(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__a21oi_1 _08461_ (.A1(_01995_),
    .A2(_02001_),
    .B1(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__a31o_1 _08462_ (.A1(_01995_),
    .A2(_02001_),
    .A3(_02005_),
    .B1(_01924_),
    .X(_02007_));
 sky130_fd_sc_hd__o221a_1 _08463_ (.A1(_01891_),
    .A2(net608),
    .B1(_02006_),
    .B2(_02007_),
    .C1(_01908_),
    .X(_00219_));
 sky130_fd_sc_hd__or3_1 _08464_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .C(_01992_),
    .X(_02008_));
 sky130_fd_sc_hd__and2_1 _08465_ (.A(_01879_),
    .B(_02008_),
    .X(_02009_));
 sky130_fd_sc_hd__xnor2_1 _08466_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _08467_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__or2_1 _08468_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02010_),
    .X(_02012_));
 sky130_fd_sc_hd__and2_1 _08469_ (.A(_02011_),
    .B(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__clkbuf_2 _08470_ (.A(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__inv_2 _08471_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ),
    .Y(_02015_));
 sky130_fd_sc_hd__o21a_1 _08472_ (.A1(_02015_),
    .A2(_02004_),
    .B1(_01995_),
    .X(_02016_));
 sky130_fd_sc_hd__a21oi_1 _08473_ (.A1(_02015_),
    .A2(_02004_),
    .B1(_02016_),
    .Y(_02017_));
 sky130_fd_sc_hd__a21o_1 _08474_ (.A1(_01998_),
    .A2(_02005_),
    .B1(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__xor2_1 _08475_ (.A(_02014_),
    .B(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _08476_ (.A0(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A1(_02019_),
    .S(_01868_),
    .X(_02020_));
 sky130_fd_sc_hd__and2_1 _08477_ (.A(_01981_),
    .B(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__clkbuf_1 _08478_ (.A(_02021_),
    .X(_00220_));
 sky130_fd_sc_hd__clkbuf_4 _08479_ (.A(_01869_),
    .X(_02022_));
 sky130_fd_sc_hd__nand2_1 _08480_ (.A(_02014_),
    .B(_02018_),
    .Y(_02023_));
 sky130_fd_sc_hd__inv_2 _08481_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ),
    .Y(_02024_));
 sky130_fd_sc_hd__inv_2 _08482_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_02025_));
 sky130_fd_sc_hd__o21a_1 _08483_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ),
    .A2(_02008_),
    .B1(_01879_),
    .X(_02026_));
 sky130_fd_sc_hd__xnor2_1 _08484_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_1 _08485_ (.A(_02024_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__nand2_1 _08486_ (.A(_02024_),
    .B(_02027_),
    .Y(_02029_));
 sky130_fd_sc_hd__and2_2 _08487_ (.A(_02028_),
    .B(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__a21oi_1 _08488_ (.A1(_02011_),
    .A2(_02023_),
    .B1(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__a31o_1 _08489_ (.A1(_02011_),
    .A2(_02023_),
    .A3(_02030_),
    .B1(_01924_),
    .X(_02032_));
 sky130_fd_sc_hd__o221a_1 _08490_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_02031_),
    .B2(_02032_),
    .C1(_01908_),
    .X(_00221_));
 sky130_fd_sc_hd__or2_1 _08491_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[8] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ),
    .X(_02033_));
 sky130_fd_sc_hd__or4_4 _08492_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .C(_01992_),
    .D(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__nand2_1 _08493_ (.A(_01880_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__xor2_1 _08494_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .B(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__nand2_1 _08495_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__or2_1 _08496_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02036_),
    .X(_02038_));
 sky130_fd_sc_hd__and2_1 _08497_ (.A(_02037_),
    .B(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__nand2_1 _08498_ (.A(_02011_),
    .B(_02028_),
    .Y(_02040_));
 sky130_fd_sc_hd__a32o_1 _08499_ (.A1(_02014_),
    .A2(_02017_),
    .A3(_02030_),
    .B1(_02040_),
    .B2(_02029_),
    .X(_02041_));
 sky130_fd_sc_hd__a41o_1 _08500_ (.A1(_01998_),
    .A2(_02005_),
    .A3(_02014_),
    .A4(_02030_),
    .B1(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__or2_1 _08501_ (.A(_02039_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__nand2_1 _08502_ (.A(_02039_),
    .B(_02042_),
    .Y(_02044_));
 sky130_fd_sc_hd__and2_1 _08503_ (.A(_02043_),
    .B(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__or2_1 _08504_ (.A(_01873_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_02046_));
 sky130_fd_sc_hd__o211a_1 _08505_ (.A1(_01867_),
    .A2(_02045_),
    .B1(_02046_),
    .C1(_01552_),
    .X(_00222_));
 sky130_fd_sc_hd__inv_2 _08506_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[10] ),
    .Y(_02047_));
 sky130_fd_sc_hd__o21a_1 _08507_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_02034_),
    .B1(_01880_),
    .X(_02048_));
 sky130_fd_sc_hd__xnor2_1 _08508_ (.A(_02047_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__and2b_1 _08509_ (.A_N(_02049_),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .X(_02050_));
 sky130_fd_sc_hd__and2b_1 _08510_ (.A_N(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .B(_02049_),
    .X(_02051_));
 sky130_fd_sc_hd__nor2_1 _08511_ (.A(_02050_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__a21oi_1 _08512_ (.A1(_02037_),
    .A2(_02044_),
    .B1(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__a31o_1 _08513_ (.A1(_02037_),
    .A2(_02044_),
    .A3(_02052_),
    .B1(_01924_),
    .X(_02054_));
 sky130_fd_sc_hd__clkbuf_4 _08514_ (.A(_01512_),
    .X(_02055_));
 sky130_fd_sc_hd__o221a_1 _08515_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_02053_),
    .B2(_02054_),
    .C1(_02055_),
    .X(_00223_));
 sky130_fd_sc_hd__or3_1 _08516_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[10] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .C(_02034_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _08517_ (.A(_01881_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__xor2_1 _08518_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__nand2_1 _08519_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__or2_1 _08520_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02058_),
    .X(_02060_));
 sky130_fd_sc_hd__and2_1 _08521_ (.A(_02059_),
    .B(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__a41oi_4 _08522_ (.A1(_01998_),
    .A2(_02005_),
    .A3(_02014_),
    .A4(_02030_),
    .B1(_02041_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(_02039_),
    .B(_02052_),
    .Y(_02063_));
 sky130_fd_sc_hd__or2b_1 _08524_ (.A(_02049_),
    .B_N(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .X(_02064_));
 sky130_fd_sc_hd__a21o_1 _08525_ (.A1(_02037_),
    .A2(_02064_),
    .B1(_02051_),
    .X(_02065_));
 sky130_fd_sc_hd__o21ai_1 _08526_ (.A1(_02062_),
    .A2(_02063_),
    .B1(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _08527_ (.A(_02061_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__o21a_1 _08528_ (.A1(_02061_),
    .A2(_02066_),
    .B1(_01868_),
    .X(_02068_));
 sky130_fd_sc_hd__a22o_1 _08529_ (.A1(_01865_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_02067_),
    .B2(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__and2_1 _08530_ (.A(_01981_),
    .B(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__clkbuf_1 _08531_ (.A(_02070_),
    .X(_00224_));
 sky130_fd_sc_hd__o21a_1 _08532_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_02056_),
    .B1(_01880_),
    .X(_02071_));
 sky130_fd_sc_hd__xor2_2 _08533_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ),
    .B(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__xnor2_2 _08534_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__a21oi_1 _08535_ (.A1(_02059_),
    .A2(_02067_),
    .B1(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__a31o_1 _08536_ (.A1(_02059_),
    .A2(_02067_),
    .A3(_02073_),
    .B1(_01924_),
    .X(_02075_));
 sky130_fd_sc_hd__o221a_1 _08537_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_02074_),
    .B2(_02075_),
    .C1(_02055_),
    .X(_00225_));
 sky130_fd_sc_hd__nand2_1 _08538_ (.A(_02061_),
    .B(_02073_),
    .Y(_02076_));
 sky130_fd_sc_hd__and2b_1 _08539_ (.A_N(_02065_),
    .B(_02073_),
    .X(_02077_));
 sky130_fd_sc_hd__inv_2 _08540_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ),
    .Y(_02078_));
 sky130_fd_sc_hd__o21a_1 _08541_ (.A1(_02078_),
    .A2(_02072_),
    .B1(_02059_),
    .X(_02079_));
 sky130_fd_sc_hd__and2_1 _08542_ (.A(_02078_),
    .B(_02072_),
    .X(_02080_));
 sky130_fd_sc_hd__o2bb2a_1 _08543_ (.A1_N(_02061_),
    .A2_N(_02077_),
    .B1(_02079_),
    .B2(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__o31a_1 _08544_ (.A1(_02062_),
    .A2(_02063_),
    .A3(_02076_),
    .B1(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__or3_1 _08545_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .C(_02056_),
    .X(_02083_));
 sky130_fd_sc_hd__and2_1 _08546_ (.A(_01881_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__xnor2_1 _08547_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .B(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _08548_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__or2_1 _08549_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02085_),
    .X(_02087_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(_02086_),
    .B(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__xor2_1 _08551_ (.A(_02082_),
    .B(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__or2_1 _08552_ (.A(_01873_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_02090_));
 sky130_fd_sc_hd__o211a_1 _08553_ (.A1(_01867_),
    .A2(_02089_),
    .B1(_02090_),
    .C1(_01552_),
    .X(_00226_));
 sky130_fd_sc_hd__inv_2 _08554_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ),
    .Y(_02091_));
 sky130_fd_sc_hd__inv_2 _08555_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[14] ),
    .Y(_02092_));
 sky130_fd_sc_hd__o21a_1 _08556_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_02083_),
    .B1(_01881_),
    .X(_02093_));
 sky130_fd_sc_hd__xnor2_2 _08557_ (.A(_02092_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__xnor2_1 _08558_ (.A(_02091_),
    .B(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__o21ai_1 _08559_ (.A1(_02082_),
    .A2(_02088_),
    .B1(_02086_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _08560_ (.A(_02095_),
    .B(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__a21o_1 _08561_ (.A1(_02095_),
    .A2(_02096_),
    .B1(_01866_),
    .X(_02098_));
 sky130_fd_sc_hd__o221a_1 _08562_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_02097_),
    .B2(_02098_),
    .C1(_02055_),
    .X(_00227_));
 sky130_fd_sc_hd__o31a_1 _08563_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[14] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .A3(_02083_),
    .B1(_01881_),
    .X(_02099_));
 sky130_fd_sc_hd__xnor2_1 _08564_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[15] ),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _08565_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__or2_1 _08566_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02100_),
    .X(_02102_));
 sky130_fd_sc_hd__and2_1 _08567_ (.A(_02101_),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__o21a_1 _08568_ (.A1(_02091_),
    .A2(_02094_),
    .B1(_02086_),
    .X(_02104_));
 sky130_fd_sc_hd__a21o_1 _08569_ (.A1(_02091_),
    .A2(_02094_),
    .B1(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__o31ai_2 _08570_ (.A1(_02082_),
    .A2(_02088_),
    .A3(_02095_),
    .B1(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(_02103_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__o21a_1 _08572_ (.A1(_02103_),
    .A2(_02106_),
    .B1(_01868_),
    .X(_02108_));
 sky130_fd_sc_hd__a22o_1 _08573_ (.A1(_01865_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_02107_),
    .B2(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__and2_1 _08574_ (.A(_01981_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__clkbuf_1 _08575_ (.A(_02110_),
    .X(_00228_));
 sky130_fd_sc_hd__or4_1 _08576_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[14] ),
    .C(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .D(_02083_),
    .X(_02111_));
 sky130_fd_sc_hd__and2_1 _08577_ (.A(_01882_),
    .B(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__xnor2_2 _08578_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__xor2_1 _08579_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ),
    .B(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__a21oi_1 _08580_ (.A1(_02101_),
    .A2(_02107_),
    .B1(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__a31o_1 _08581_ (.A1(_02101_),
    .A2(_02107_),
    .A3(_02114_),
    .B1(_01924_),
    .X(_02116_));
 sky130_fd_sc_hd__o221a_1 _08582_ (.A1(_02022_),
    .A2(net499),
    .B1(_02115_),
    .B2(_02116_),
    .C1(_02055_),
    .X(_00229_));
 sky130_fd_sc_hd__inv_2 _08583_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _08584_ (.A(_01877_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__a21bo_1 _08585_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_02113_),
    .B1_N(_02101_),
    .X(_02119_));
 sky130_fd_sc_hd__o21ai_1 _08586_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_02113_),
    .B1(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand3_1 _08587_ (.A(_02103_),
    .B(_02106_),
    .C(_02114_),
    .Y(_02121_));
 sky130_fd_sc_hd__nor2_1 _08588_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02111_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _08589_ (.A(_01549_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__mux2_1 _08590_ (.A0(_02123_),
    .A1(_01549_),
    .S(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[17] ),
    .X(_02124_));
 sky130_fd_sc_hd__a21oi_1 _08591_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_02122_),
    .B1(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__and2_1 _08592_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__nor2_1 _08593_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02125_),
    .Y(_02127_));
 sky130_fd_sc_hd__or2_1 _08594_ (.A(_02126_),
    .B(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__a21oi_1 _08595_ (.A1(_02120_),
    .A2(_02121_),
    .B1(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__a31o_1 _08596_ (.A1(_02128_),
    .A2(_02120_),
    .A3(_02121_),
    .B1(_01865_),
    .X(_02130_));
 sky130_fd_sc_hd__nor2_1 _08597_ (.A(_02129_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__clkbuf_8 _08598_ (.A(_01794_),
    .X(_02132_));
 sky130_fd_sc_hd__o21a_1 _08599_ (.A1(_02118_),
    .A2(_02131_),
    .B1(_02132_),
    .X(_00230_));
 sky130_fd_sc_hd__xor2_1 _08600_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[17] ),
    .B(_02124_),
    .X(_02133_));
 sky130_fd_sc_hd__o21a_1 _08601_ (.A1(_02126_),
    .A2(_02129_),
    .B1(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__o31ai_1 _08602_ (.A1(_02126_),
    .A2(_02129_),
    .A3(_02133_),
    .B1(_01870_),
    .Y(_02135_));
 sky130_fd_sc_hd__o221a_1 _08603_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B1(_02134_),
    .B2(_02135_),
    .C1(_02055_),
    .X(_00231_));
 sky130_fd_sc_hd__and2_1 _08604_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ),
    .X(_02136_));
 sky130_fd_sc_hd__nor2_1 _08605_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ),
    .Y(_02137_));
 sky130_fd_sc_hd__o21ai_1 _08606_ (.A1(_02136_),
    .A2(_02137_),
    .B1(_01877_),
    .Y(_02138_));
 sky130_fd_sc_hd__o211a_1 _08607_ (.A1(_01876_),
    .A2(net273),
    .B1(_01945_),
    .C1(_02138_),
    .X(_00232_));
 sky130_fd_sc_hd__and2b_1 _08608_ (.A_N(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .X(_02139_));
 sky130_fd_sc_hd__xnor2_1 _08609_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__xnor2_1 _08610_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nor2_1 _08611_ (.A(_02136_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__and2_1 _08612_ (.A(_02136_),
    .B(_02141_),
    .X(_02143_));
 sky130_fd_sc_hd__o21ai_1 _08613_ (.A1(_02142_),
    .A2(_02143_),
    .B1(_01877_),
    .Y(_02144_));
 sky130_fd_sc_hd__o211a_1 _08614_ (.A1(_01876_),
    .A2(net310),
    .B1(_01945_),
    .C1(_02144_),
    .X(_00233_));
 sky130_fd_sc_hd__nor2_1 _08615_ (.A(_01961_),
    .B(_02140_),
    .Y(_02145_));
 sky130_fd_sc_hd__inv_2 _08616_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_02146_));
 sky130_fd_sc_hd__o21a_1 _08617_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B1(_01879_),
    .X(_02147_));
 sky130_fd_sc_hd__xnor2_1 _08618_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__xnor2_1 _08619_ (.A(_02146_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__o21bai_2 _08620_ (.A1(_02145_),
    .A2(_02143_),
    .B1_N(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__or3b_1 _08621_ (.A(_02145_),
    .B(_02143_),
    .C_N(_02149_),
    .X(_02151_));
 sky130_fd_sc_hd__inv_2 _08622_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_02152_));
 sky130_fd_sc_hd__nor2_1 _08623_ (.A(_01868_),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__a31o_1 _08624_ (.A1(_01869_),
    .A2(_02150_),
    .A3(_02151_),
    .B1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__and2_1 _08625_ (.A(_01981_),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__clkbuf_1 _08626_ (.A(_02155_),
    .X(_00234_));
 sky130_fd_sc_hd__inv_2 _08627_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_02156_));
 sky130_fd_sc_hd__or2_1 _08628_ (.A(_02146_),
    .B(_02148_),
    .X(_02157_));
 sky130_fd_sc_hd__inv_2 _08629_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_02158_));
 sky130_fd_sc_hd__o31a_1 _08630_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .A3(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .B1(_01879_),
    .X(_02159_));
 sky130_fd_sc_hd__xnor2_1 _08631_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ),
    .B(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hd__nor2_1 _08632_ (.A(_02158_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__and2_1 _08633_ (.A(_02158_),
    .B(_02160_),
    .X(_02162_));
 sky130_fd_sc_hd__or2_1 _08634_ (.A(_02161_),
    .B(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__and3_1 _08635_ (.A(_02157_),
    .B(_02150_),
    .C(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__a21oi_2 _08636_ (.A1(_02157_),
    .A2(_02150_),
    .B1(_02163_),
    .Y(_02165_));
 sky130_fd_sc_hd__or3_1 _08637_ (.A(_01864_),
    .B(_02164_),
    .C(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__o21a_1 _08638_ (.A1(_01869_),
    .A2(_02156_),
    .B1(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__and2b_1 _08639_ (.A_N(_02167_),
    .B(_01979_),
    .X(_02168_));
 sky130_fd_sc_hd__clkbuf_1 _08640_ (.A(_02168_),
    .X(_00235_));
 sky130_fd_sc_hd__inv_2 _08641_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_02169_));
 sky130_fd_sc_hd__or4_4 _08642_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ),
    .C(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .D(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ),
    .X(_02170_));
 sky130_fd_sc_hd__nand2_1 _08643_ (.A(_01879_),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__xnor2_1 _08644_ (.A(_02015_),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor2_1 _08645_ (.A(_02169_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__and2_1 _08646_ (.A(_02169_),
    .B(_02172_),
    .X(_02174_));
 sky130_fd_sc_hd__or2_1 _08647_ (.A(_02173_),
    .B(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__inv_2 _08648_ (.A(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__o21a_1 _08649_ (.A1(_02161_),
    .A2(_02165_),
    .B1(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__or3_1 _08650_ (.A(_02161_),
    .B(_02165_),
    .C(_02176_),
    .X(_02178_));
 sky130_fd_sc_hd__and2b_1 _08651_ (.A_N(_02177_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__or2_1 _08652_ (.A(_01873_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_02180_));
 sky130_fd_sc_hd__o211a_1 _08653_ (.A1(_01867_),
    .A2(_02179_),
    .B1(_02180_),
    .C1(_01552_),
    .X(_00236_));
 sky130_fd_sc_hd__o21a_1 _08654_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_02170_),
    .B1(_01879_),
    .X(_02181_));
 sky130_fd_sc_hd__xor2_1 _08655_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__and2_1 _08656_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .B(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__or2_1 _08657_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ),
    .B(_02182_),
    .X(_02184_));
 sky130_fd_sc_hd__and2b_1 _08658_ (.A_N(_02183_),
    .B(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__nor2_1 _08659_ (.A(_02173_),
    .B(_02177_),
    .Y(_02186_));
 sky130_fd_sc_hd__xnor2_1 _08660_ (.A(_02185_),
    .B(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__or2_1 _08661_ (.A(_01873_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_02188_));
 sky130_fd_sc_hd__o211a_1 _08662_ (.A1(_01866_),
    .A2(_02187_),
    .B1(_02188_),
    .C1(_01552_),
    .X(_00237_));
 sky130_fd_sc_hd__and2_1 _08663_ (.A(_02177_),
    .B(_02185_),
    .X(_02189_));
 sky130_fd_sc_hd__o21a_1 _08664_ (.A1(_02173_),
    .A2(_02183_),
    .B1(_02184_),
    .X(_02190_));
 sky130_fd_sc_hd__or3_1 _08665_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ),
    .C(_02170_),
    .X(_02191_));
 sky130_fd_sc_hd__and2_1 _08666_ (.A(_01880_),
    .B(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__xnor2_2 _08667_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__xnor2_2 _08668_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__o21ai_1 _08669_ (.A1(_02189_),
    .A2(_02190_),
    .B1(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__o31a_1 _08670_ (.A1(_02194_),
    .A2(_02189_),
    .A3(_02190_),
    .B1(_01868_),
    .X(_02196_));
 sky130_fd_sc_hd__a22o_1 _08671_ (.A1(_01865_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1(_02195_),
    .B2(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__and2_1 _08672_ (.A(_01981_),
    .B(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__clkbuf_1 _08673_ (.A(_02198_),
    .X(_00238_));
 sky130_fd_sc_hd__or2_1 _08674_ (.A(_02002_),
    .B(_02193_),
    .X(_02199_));
 sky130_fd_sc_hd__o21a_1 _08675_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ),
    .A2(_02191_),
    .B1(_01879_),
    .X(_02200_));
 sky130_fd_sc_hd__xor2_1 _08676_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__nand2_1 _08677_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__or2_1 _08678_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02201_),
    .X(_02203_));
 sky130_fd_sc_hd__and2_1 _08679_ (.A(_02202_),
    .B(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__a21oi_1 _08680_ (.A1(_02199_),
    .A2(_02195_),
    .B1(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__a31o_1 _08681_ (.A1(_02199_),
    .A2(_02195_),
    .A3(_02204_),
    .B1(_01924_),
    .X(_02206_));
 sky130_fd_sc_hd__o221a_1 _08682_ (.A1(_02022_),
    .A2(net574),
    .B1(_02205_),
    .B2(_02206_),
    .C1(_02055_),
    .X(_00239_));
 sky130_fd_sc_hd__or2_1 _08683_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ),
    .X(_02207_));
 sky130_fd_sc_hd__or4_4 _08684_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ),
    .C(_02170_),
    .D(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__nand2_1 _08685_ (.A(_01880_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__xor2_1 _08686_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .B(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__or2_1 _08687_ (.A(_02025_),
    .B(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(_02025_),
    .B(_02210_),
    .Y(_02212_));
 sky130_fd_sc_hd__nand2_1 _08689_ (.A(_02211_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__o2111a_1 _08690_ (.A1(_02161_),
    .A2(_02165_),
    .B1(_02176_),
    .C1(_02185_),
    .D1(_02204_),
    .X(_02214_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(_02199_),
    .B(_02202_),
    .Y(_02215_));
 sky130_fd_sc_hd__a32o_1 _08692_ (.A1(_02194_),
    .A2(_02190_),
    .A3(_02204_),
    .B1(_02215_),
    .B2(_02203_),
    .X(_02216_));
 sky130_fd_sc_hd__a21o_1 _08693_ (.A1(_02194_),
    .A2(_02214_),
    .B1(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__xnor2_1 _08694_ (.A(_02213_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__or2_1 _08695_ (.A(_01873_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_02219_));
 sky130_fd_sc_hd__o211a_1 _08696_ (.A1(_01866_),
    .A2(_02218_),
    .B1(_02219_),
    .C1(_01552_),
    .X(_00240_));
 sky130_fd_sc_hd__o21a_1 _08697_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_02208_),
    .B1(_01880_),
    .X(_02220_));
 sky130_fd_sc_hd__xor2_2 _08698_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__xnor2_1 _08699_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__a21oi_1 _08700_ (.A1(_02194_),
    .A2(_02214_),
    .B1(_02216_),
    .Y(_02223_));
 sky130_fd_sc_hd__o21ai_1 _08701_ (.A1(_02213_),
    .A2(_02223_),
    .B1(_02211_),
    .Y(_02224_));
 sky130_fd_sc_hd__nor2_1 _08702_ (.A(_02222_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__a21o_1 _08703_ (.A1(_02222_),
    .A2(_02224_),
    .B1(_01866_),
    .X(_02226_));
 sky130_fd_sc_hd__o221a_1 _08704_ (.A1(_02022_),
    .A2(net581),
    .B1(_02225_),
    .B2(_02226_),
    .C1(_02055_),
    .X(_00241_));
 sky130_fd_sc_hd__a21bo_1 _08705_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_02221_),
    .B1_N(_02211_),
    .X(_02227_));
 sky130_fd_sc_hd__o21a_1 _08706_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_02221_),
    .B1(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__inv_2 _08707_ (.A(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__or3_1 _08708_ (.A(_02213_),
    .B(_02223_),
    .C(_02222_),
    .X(_02230_));
 sky130_fd_sc_hd__or3_1 _08709_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ),
    .C(_02208_),
    .X(_02231_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_01881_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__xor2_1 _08711_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ),
    .B(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__xnor2_1 _08712_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[10] ),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__a21bo_1 _08713_ (.A1(_02229_),
    .A2(_02230_),
    .B1_N(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__or3b_1 _08714_ (.A(_02234_),
    .B(_02228_),
    .C_N(_02230_),
    .X(_02236_));
 sky130_fd_sc_hd__inv_2 _08715_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .Y(_02237_));
 sky130_fd_sc_hd__nor2_1 _08716_ (.A(_01868_),
    .B(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__a31o_1 _08717_ (.A1(_01869_),
    .A2(_02235_),
    .A3(_02236_),
    .B1(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__and2_1 _08718_ (.A(_01981_),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_1 _08719_ (.A(_02240_),
    .X(_00242_));
 sky130_fd_sc_hd__or2_1 _08720_ (.A(_02047_),
    .B(_02233_),
    .X(_02241_));
 sky130_fd_sc_hd__o21a_1 _08721_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_02231_),
    .B1(_01880_),
    .X(_02242_));
 sky130_fd_sc_hd__xor2_1 _08722_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__and2_1 _08723_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__nor2_1 _08724_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02243_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _08725_ (.A(_02244_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21oi_1 _08726_ (.A1(_02241_),
    .A2(_02235_),
    .B1(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__a31o_1 _08727_ (.A1(_02241_),
    .A2(_02235_),
    .A3(_02246_),
    .B1(_01865_),
    .X(_02248_));
 sky130_fd_sc_hd__o221a_1 _08728_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_02247_),
    .B2(_02248_),
    .C1(_02055_),
    .X(_00243_));
 sky130_fd_sc_hd__or3_2 _08729_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ),
    .C(_02231_),
    .X(_02249_));
 sky130_fd_sc_hd__and2_1 _08730_ (.A(_01881_),
    .B(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__xnor2_2 _08731_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__xor2_2 _08732_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ),
    .B(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__and4bb_1 _08733_ (.A_N(_02213_),
    .B_N(_02222_),
    .C(_02234_),
    .D(_02246_),
    .X(_02253_));
 sky130_fd_sc_hd__and3_1 _08734_ (.A(_02234_),
    .B(_02228_),
    .C(_02246_),
    .X(_02254_));
 sky130_fd_sc_hd__nand2_1 _08735_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02243_),
    .Y(_02255_));
 sky130_fd_sc_hd__a21oi_1 _08736_ (.A1(_02241_),
    .A2(_02255_),
    .B1(_02245_),
    .Y(_02256_));
 sky130_fd_sc_hd__a211o_1 _08737_ (.A1(_02217_),
    .A2(_02253_),
    .B1(_02254_),
    .C1(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__xnor2_1 _08738_ (.A(_02252_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__or2_1 _08739_ (.A(_01869_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_02259_));
 sky130_fd_sc_hd__buf_4 _08740_ (.A(_01474_),
    .X(_02260_));
 sky130_fd_sc_hd__o211a_1 _08741_ (.A1(_01866_),
    .A2(_02258_),
    .B1(_02259_),
    .C1(_02260_),
    .X(_00244_));
 sky130_fd_sc_hd__o21a_1 _08742_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_02249_),
    .B1(_01881_),
    .X(_02261_));
 sky130_fd_sc_hd__xor2_2 _08743_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__xnor2_1 _08744_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__inv_2 _08745_ (.A(_02251_),
    .Y(_02264_));
 sky130_fd_sc_hd__and2b_1 _08746_ (.A_N(_02252_),
    .B(_02257_),
    .X(_02265_));
 sky130_fd_sc_hd__a21o_1 _08747_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_02264_),
    .B1(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__nor2_1 _08748_ (.A(_02263_),
    .B(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21o_1 _08749_ (.A1(_02263_),
    .A2(_02266_),
    .B1(_01866_),
    .X(_02268_));
 sky130_fd_sc_hd__o221a_1 _08750_ (.A1(_02022_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_02267_),
    .B2(_02268_),
    .C1(_02055_),
    .X(_00245_));
 sky130_fd_sc_hd__a22o_1 _08751_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_02264_),
    .B1(_02262_),
    .B2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .X(_02269_));
 sky130_fd_sc_hd__o21ai_2 _08752_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_02262_),
    .B1(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _08753_ (.A(_02252_),
    .B(_02263_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(_02257_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__o31a_1 _08755_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ),
    .A2(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ),
    .A3(_02249_),
    .B1(_01881_),
    .X(_02273_));
 sky130_fd_sc_hd__xnor2_1 _08756_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__or2_1 _08757_ (.A(_02092_),
    .B(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__nand2_1 _08758_ (.A(_02092_),
    .B(_02274_),
    .Y(_02276_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(_02275_),
    .B(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__a21o_1 _08760_ (.A1(_02270_),
    .A2(_02272_),
    .B1(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__a31oi_1 _08761_ (.A1(_02277_),
    .A2(_02270_),
    .A3(_02272_),
    .B1(_01865_),
    .Y(_02279_));
 sky130_fd_sc_hd__a22o_1 _08762_ (.A1(_01865_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_02278_),
    .B2(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__and2_1 _08763_ (.A(_01981_),
    .B(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__clkbuf_1 _08764_ (.A(_02281_),
    .X(_00246_));
 sky130_fd_sc_hd__inv_2 _08765_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[15] ),
    .Y(_02282_));
 sky130_fd_sc_hd__or4_4 _08766_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ),
    .C(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ),
    .D(_02249_),
    .X(_02283_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(_01881_),
    .B(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__xor2_2 _08768_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__xnor2_1 _08769_ (.A(_02282_),
    .B(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_1 _08770_ (.A(_02275_),
    .B(_02278_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _08771_ (.A(_02286_),
    .B(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__a21o_1 _08772_ (.A1(_02286_),
    .A2(_02287_),
    .B1(_01924_),
    .X(_02289_));
 sky130_fd_sc_hd__o221a_1 _08773_ (.A1(_01877_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_02288_),
    .B2(_02289_),
    .C1(_02055_),
    .X(_00247_));
 sky130_fd_sc_hd__and2_1 _08774_ (.A(_01924_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .X(_02290_));
 sky130_fd_sc_hd__nor2_1 _08775_ (.A(_02277_),
    .B(_02286_),
    .Y(_02291_));
 sky130_fd_sc_hd__and3_1 _08776_ (.A(_02257_),
    .B(_02271_),
    .C(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__o21a_1 _08777_ (.A1(_02282_),
    .A2(_02285_),
    .B1(_02275_),
    .X(_02293_));
 sky130_fd_sc_hd__a21oi_1 _08778_ (.A1(_02282_),
    .A2(_02285_),
    .B1(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__and2b_1 _08779_ (.A_N(_02270_),
    .B(_02291_),
    .X(_02295_));
 sky130_fd_sc_hd__nor2_2 _08780_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02283_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _08781_ (.A(_01549_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__mux2_1 _08782_ (.A0(_02297_),
    .A1(_01549_),
    .S(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[17] ),
    .X(_02298_));
 sky130_fd_sc_hd__a21o_1 _08783_ (.A1(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[17] ),
    .A2(_02296_),
    .B1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__xor2_1 _08784_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__o31a_1 _08785_ (.A1(_02292_),
    .A2(_02294_),
    .A3(_02295_),
    .B1(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__or4_1 _08786_ (.A(_02300_),
    .B(_02292_),
    .C(_02294_),
    .D(_02295_),
    .X(_02302_));
 sky130_fd_sc_hd__and3b_1 _08787_ (.A_N(_02301_),
    .B(_02302_),
    .C(_01873_),
    .X(_02303_));
 sky130_fd_sc_hd__o21a_1 _08788_ (.A1(_02290_),
    .A2(_02303_),
    .B1(_02132_),
    .X(_00248_));
 sky130_fd_sc_hd__and2_1 _08789_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02299_),
    .X(_02304_));
 sky130_fd_sc_hd__xnor2_1 _08790_ (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[17] ),
    .B(_02298_),
    .Y(_02305_));
 sky130_fd_sc_hd__o21a_1 _08791_ (.A1(_02304_),
    .A2(_02301_),
    .B1(_02305_),
    .X(_02306_));
 sky130_fd_sc_hd__o31ai_1 _08792_ (.A1(_02304_),
    .A2(_02301_),
    .A3(_02305_),
    .B1(_01870_),
    .Y(_02307_));
 sky130_fd_sc_hd__clkbuf_4 _08793_ (.A(_01252_),
    .X(_02308_));
 sky130_fd_sc_hd__clkbuf_4 _08794_ (.A(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__o221a_1 _08795_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_01876_),
    .B1(_02306_),
    .B2(_02307_),
    .C1(_02309_),
    .X(_00249_));
 sky130_fd_sc_hd__buf_4 _08796_ (.A(_01252_),
    .X(_02310_));
 sky130_fd_sc_hd__and2_1 _08797_ (.A(_01870_),
    .B(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__clkbuf_1 _08798_ (.A(_02311_),
    .X(_00250_));
 sky130_fd_sc_hd__inv_2 _08799_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_02312_));
 sky130_fd_sc_hd__clkbuf_4 _08800_ (.A(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__buf_4 _08801_ (.A(_02313_),
    .X(_02314_));
 sky130_fd_sc_hd__clkbuf_4 _08802_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02315_));
 sky130_fd_sc_hd__or2_1 _08803_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_02315_),
    .X(_02316_));
 sky130_fd_sc_hd__o211a_1 _08804_ (.A1(_02314_),
    .A2(net155),
    .B1(_01945_),
    .C1(_02316_),
    .X(_00251_));
 sky130_fd_sc_hd__or2_1 _08805_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_02315_),
    .X(_02317_));
 sky130_fd_sc_hd__o211a_1 _08806_ (.A1(_02314_),
    .A2(net191),
    .B1(_01945_),
    .C1(_02317_),
    .X(_00252_));
 sky130_fd_sc_hd__or2_1 _08807_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_02318_));
 sky130_fd_sc_hd__o211a_1 _08808_ (.A1(_02314_),
    .A2(net147),
    .B1(_01945_),
    .C1(_02318_),
    .X(_00253_));
 sky130_fd_sc_hd__clkbuf_4 _08809_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02319_));
 sky130_fd_sc_hd__clkbuf_4 _08810_ (.A(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__clkbuf_4 _08811_ (.A(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__buf_4 _08812_ (.A(_02319_),
    .X(_02322_));
 sky130_fd_sc_hd__nand2_1 _08813_ (.A(_02322_),
    .B(net300),
    .Y(_02323_));
 sky130_fd_sc_hd__o211a_1 _08814_ (.A1(_02321_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B1(_01945_),
    .C1(_02323_),
    .X(_00254_));
 sky130_fd_sc_hd__or2_1 _08815_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(_02324_));
 sky130_fd_sc_hd__nand2_1 _08816_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .Y(_02325_));
 sky130_fd_sc_hd__and3_1 _08817_ (.A(_01959_),
    .B(_02324_),
    .C(_02325_),
    .X(_02326_));
 sky130_fd_sc_hd__a21oi_1 _08818_ (.A1(_02324_),
    .A2(_02325_),
    .B1(_01959_),
    .Y(_02327_));
 sky130_fd_sc_hd__o21ai_1 _08819_ (.A1(_02326_),
    .A2(_02327_),
    .B1(_02322_),
    .Y(_02328_));
 sky130_fd_sc_hd__o211a_1 _08820_ (.A1(_02321_),
    .A2(net364),
    .B1(_01945_),
    .C1(_02328_),
    .X(_00255_));
 sky130_fd_sc_hd__clkbuf_4 _08821_ (.A(_02315_),
    .X(_02329_));
 sky130_fd_sc_hd__or2_1 _08822_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_02324_),
    .X(_02330_));
 sky130_fd_sc_hd__nand2_1 _08823_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_02324_),
    .Y(_02331_));
 sky130_fd_sc_hd__a21oi_1 _08824_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_02327_),
    .Y(_02332_));
 sky130_fd_sc_hd__buf_4 _08825_ (.A(_02312_),
    .X(_02333_));
 sky130_fd_sc_hd__a31o_1 _08826_ (.A1(_02327_),
    .A2(_02330_),
    .A3(_02331_),
    .B1(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__o221a_1 _08827_ (.A1(_02329_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B1(_02332_),
    .B2(_02334_),
    .C1(_02309_),
    .X(_00256_));
 sky130_fd_sc_hd__and3_1 _08828_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .C(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(_02335_));
 sky130_fd_sc_hd__or2_1 _08829_ (.A(_01958_),
    .B(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_1 _08830_ (.A(_01958_),
    .B(_02330_),
    .Y(_02337_));
 sky130_fd_sc_hd__a21oi_1 _08831_ (.A1(_02336_),
    .A2(_02337_),
    .B1(net588),
    .Y(_02338_));
 sky130_fd_sc_hd__a31o_1 _08832_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_02336_),
    .A3(_02337_),
    .B1(_02333_),
    .X(_02339_));
 sky130_fd_sc_hd__o221a_1 _08833_ (.A1(_02329_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B1(_02338_),
    .B2(_02339_),
    .C1(_02309_),
    .X(_00257_));
 sky130_fd_sc_hd__o21ai_1 _08834_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_02335_),
    .B1(_02337_),
    .Y(_02340_));
 sky130_fd_sc_hd__inv_2 _08835_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_02341_));
 sky130_fd_sc_hd__buf_2 _08836_ (.A(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__buf_2 _08837_ (.A(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__clkbuf_4 _08838_ (.A(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__or2_1 _08839_ (.A(_02344_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(_02345_));
 sky130_fd_sc_hd__a21oi_1 _08840_ (.A1(_02340_),
    .A2(_02345_),
    .B1(net469),
    .Y(_02346_));
 sky130_fd_sc_hd__a31o_1 _08841_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(_02340_),
    .A3(_02345_),
    .B1(_02333_),
    .X(_02347_));
 sky130_fd_sc_hd__o221a_1 _08842_ (.A1(_02329_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B1(_02346_),
    .B2(_02347_),
    .C1(_02309_),
    .X(_00258_));
 sky130_fd_sc_hd__a21o_1 _08843_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_02330_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(_02348_));
 sky130_fd_sc_hd__o21a_1 _08844_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_02335_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(_02349_));
 sky130_fd_sc_hd__inv_2 _08845_ (.A(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__mux2_1 _08846_ (.A0(_02348_),
    .A1(_02350_),
    .S(_02344_),
    .X(_02351_));
 sky130_fd_sc_hd__xnor2_1 _08847_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(_02322_),
    .B(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__o211a_1 _08849_ (.A1(_02321_),
    .A2(net355),
    .B1(_01945_),
    .C1(_02353_),
    .X(_00259_));
 sky130_fd_sc_hd__a21oi_1 _08850_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_02348_),
    .B1(_02344_),
    .Y(_02354_));
 sky130_fd_sc_hd__o21a_1 _08851_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_02349_),
    .B1(_02344_),
    .X(_02355_));
 sky130_fd_sc_hd__inv_2 _08852_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_02356_));
 sky130_fd_sc_hd__o21a_1 _08853_ (.A1(_02354_),
    .A2(_02355_),
    .B1(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__o31ai_1 _08854_ (.A1(_02356_),
    .A2(_02354_),
    .A3(_02355_),
    .B1(_02320_),
    .Y(_02358_));
 sky130_fd_sc_hd__o221a_1 _08855_ (.A1(_02329_),
    .A2(net582),
    .B1(_02357_),
    .B2(_02358_),
    .C1(_02309_),
    .X(_00260_));
 sky130_fd_sc_hd__a21oi_1 _08856_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_02348_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_02359_));
 sky130_fd_sc_hd__o22a_1 _08857_ (.A1(_01959_),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B1(_02355_),
    .B2(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__xor2_1 _08858_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__or2_1 _08859_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(_02362_));
 sky130_fd_sc_hd__o211a_1 _08860_ (.A1(_02314_),
    .A2(_02361_),
    .B1(_02362_),
    .C1(_02260_),
    .X(_00261_));
 sky130_fd_sc_hd__or2b_1 _08861_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B_N(_02359_),
    .X(_02363_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(_01959_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__o211a_1 _08863_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_02349_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(_02365_));
 sky130_fd_sc_hd__or2_1 _08864_ (.A(_01958_),
    .B(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__inv_2 _08865_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_02367_));
 sky130_fd_sc_hd__a21oi_1 _08866_ (.A1(_02364_),
    .A2(_02366_),
    .B1(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__buf_4 _08867_ (.A(_02313_),
    .X(_02369_));
 sky130_fd_sc_hd__a31o_1 _08868_ (.A1(_02367_),
    .A2(_02364_),
    .A3(_02366_),
    .B1(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__o221a_1 _08869_ (.A1(_02329_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_02368_),
    .B2(_02370_),
    .C1(_02309_),
    .X(_00262_));
 sky130_fd_sc_hd__or2_1 _08870_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_02363_),
    .X(_02371_));
 sky130_fd_sc_hd__nand2_1 _08871_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_02365_),
    .Y(_02372_));
 sky130_fd_sc_hd__mux2_1 _08872_ (.A0(_02371_),
    .A1(_02372_),
    .S(_02344_),
    .X(_02373_));
 sky130_fd_sc_hd__and2_1 _08873_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__o21ai_1 _08874_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_02373_),
    .B1(_02320_),
    .Y(_02375_));
 sky130_fd_sc_hd__o221a_1 _08875_ (.A1(_02329_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_02374_),
    .B2(_02375_),
    .C1(_02309_),
    .X(_00263_));
 sky130_fd_sc_hd__and3_1 _08876_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(_02365_),
    .X(_02376_));
 sky130_fd_sc_hd__o21ai_1 _08877_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_02371_),
    .B1(_01959_),
    .Y(_02377_));
 sky130_fd_sc_hd__o21ai_1 _08878_ (.A1(_01959_),
    .A2(_02376_),
    .B1(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__xnor2_1 _08879_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__or2_1 _08880_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(_02380_));
 sky130_fd_sc_hd__o211a_1 _08881_ (.A1(_02314_),
    .A2(_02379_),
    .B1(_02380_),
    .C1(_02260_),
    .X(_00264_));
 sky130_fd_sc_hd__clkbuf_4 _08882_ (.A(_01455_),
    .X(_02381_));
 sky130_fd_sc_hd__a21oi_1 _08883_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_02376_),
    .B1(_01958_),
    .Y(_02382_));
 sky130_fd_sc_hd__or3_1 _08884_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_02371_),
    .X(_02383_));
 sky130_fd_sc_hd__a21bo_1 _08885_ (.A1(_01959_),
    .A2(_02383_),
    .B1_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(_02384_));
 sky130_fd_sc_hd__a21oi_1 _08886_ (.A1(_01959_),
    .A2(_02383_),
    .B1(_02382_),
    .Y(_02385_));
 sky130_fd_sc_hd__o221ai_1 _08887_ (.A1(_02382_),
    .A2(_02384_),
    .B1(_02385_),
    .B2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C1(_02320_),
    .Y(_02386_));
 sky130_fd_sc_hd__o211a_1 _08888_ (.A1(_02321_),
    .A2(net447),
    .B1(_02381_),
    .C1(_02386_),
    .X(_00265_));
 sky130_fd_sc_hd__clkbuf_4 _08889_ (.A(_02319_),
    .X(_02387_));
 sky130_fd_sc_hd__or2_1 _08890_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_02382_),
    .X(_02388_));
 sky130_fd_sc_hd__inv_2 _08891_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .Y(_02389_));
 sky130_fd_sc_hd__a21oi_1 _08892_ (.A1(_02384_),
    .A2(_02388_),
    .B1(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__a31o_1 _08893_ (.A1(_02389_),
    .A2(_02384_),
    .A3(_02388_),
    .B1(_02369_),
    .X(_02391_));
 sky130_fd_sc_hd__o221a_1 _08894_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_02390_),
    .B2(_02391_),
    .C1(_02309_),
    .X(_00266_));
 sky130_fd_sc_hd__inv_2 _08895_ (.A(net481),
    .Y(_02392_));
 sky130_fd_sc_hd__and3_1 _08896_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C(_02383_),
    .X(_02393_));
 sky130_fd_sc_hd__a211o_1 _08897_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_02376_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(_02394_));
 sky130_fd_sc_hd__inv_2 _08898_ (.A(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(_02393_),
    .A1(_02395_),
    .S(_02344_),
    .X(_02396_));
 sky130_fd_sc_hd__a21oi_1 _08900_ (.A1(_02392_),
    .A2(_02396_),
    .B1(_02333_),
    .Y(_02397_));
 sky130_fd_sc_hd__o21ai_1 _08901_ (.A1(_02392_),
    .A2(_02396_),
    .B1(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__o211a_1 _08902_ (.A1(_02321_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_02381_),
    .C1(_02398_),
    .X(_00267_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_02394_),
    .X(_02399_));
 sky130_fd_sc_hd__and3_1 _08904_ (.A(_01958_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .C(_02393_),
    .X(_02400_));
 sky130_fd_sc_hd__o21ba_1 _08905_ (.A1(_01959_),
    .A2(_02399_),
    .B1_N(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__and2_1 _08906_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__o21ai_1 _08907_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_02401_),
    .B1(_02320_),
    .Y(_02403_));
 sky130_fd_sc_hd__o221a_1 _08908_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_02402_),
    .B2(_02403_),
    .C1(_02309_),
    .X(_00268_));
 sky130_fd_sc_hd__o21ai_1 _08909_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_02399_),
    .B1(_02344_),
    .Y(_02404_));
 sky130_fd_sc_hd__a31o_1 _08910_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_02393_),
    .B1(_02344_),
    .X(_02405_));
 sky130_fd_sc_hd__inv_2 _08911_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .Y(_02406_));
 sky130_fd_sc_hd__a21oi_1 _08912_ (.A1(_02404_),
    .A2(_02405_),
    .B1(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__a31o_1 _08913_ (.A1(_02406_),
    .A2(_02404_),
    .A3(_02405_),
    .B1(_02369_),
    .X(_02408_));
 sky130_fd_sc_hd__o221a_1 _08914_ (.A1(_02387_),
    .A2(net440),
    .B1(_02407_),
    .B2(_02408_),
    .C1(_02309_),
    .X(_00269_));
 sky130_fd_sc_hd__clkbuf_4 _08915_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_02409_));
 sky130_fd_sc_hd__nand2_1 _08916_ (.A(net531),
    .B(_02405_),
    .Y(_02410_));
 sky130_fd_sc_hd__a21o_1 _08917_ (.A1(_02404_),
    .A2(_02410_),
    .B1(_02314_),
    .X(_02411_));
 sky130_fd_sc_hd__o211a_1 _08918_ (.A1(_02321_),
    .A2(_02409_),
    .B1(_02381_),
    .C1(_02411_),
    .X(_00270_));
 sky130_fd_sc_hd__nor2_1 _08919_ (.A(_02152_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_02412_));
 sky130_fd_sc_hd__a21o_1 _08920_ (.A1(_02152_),
    .A2(net649),
    .B1(_02333_),
    .X(_02413_));
 sky130_fd_sc_hd__clkbuf_4 _08921_ (.A(_02308_),
    .X(_02414_));
 sky130_fd_sc_hd__o221a_1 _08922_ (.A1(_02387_),
    .A2(net449),
    .B1(_02412_),
    .B2(_02413_),
    .C1(_02414_),
    .X(_00271_));
 sky130_fd_sc_hd__and2b_1 _08923_ (.A_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__xnor2_1 _08924_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__xnor2_1 _08925_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__xor2_1 _08926_ (.A(_02412_),
    .B(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__or2_1 _08927_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_02419_));
 sky130_fd_sc_hd__o211a_1 _08928_ (.A1(_02314_),
    .A2(_02418_),
    .B1(_02419_),
    .C1(_02260_),
    .X(_00272_));
 sky130_fd_sc_hd__and2_1 _08929_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_02416_),
    .X(_02420_));
 sky130_fd_sc_hd__nor2_1 _08930_ (.A(_02412_),
    .B(_02417_),
    .Y(_02421_));
 sky130_fd_sc_hd__o21ba_1 _08931_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_02422_));
 sky130_fd_sc_hd__xnor2_1 _08932_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__nand2_1 _08933_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__or2_1 _08934_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_02423_),
    .X(_02425_));
 sky130_fd_sc_hd__and2_1 _08935_ (.A(_02424_),
    .B(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__o21ai_2 _08936_ (.A1(_02420_),
    .A2(_02421_),
    .B1(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__o31a_1 _08937_ (.A1(_02420_),
    .A2(_02421_),
    .A3(_02426_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02428_));
 sky130_fd_sc_hd__a22oi_1 _08938_ (.A1(_02313_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_02427_),
    .B2(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__and2b_1 _08939_ (.A_N(_02429_),
    .B(_01979_),
    .X(_02430_));
 sky130_fd_sc_hd__clkbuf_1 _08940_ (.A(_02430_),
    .X(_00273_));
 sky130_fd_sc_hd__o31a_1 _08941_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A3(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_02341_),
    .X(_02431_));
 sky130_fd_sc_hd__xnor2_1 _08942_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__and2_1 _08943_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__nor2_1 _08944_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_02432_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _08945_ (.A(_02433_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__nand2_1 _08946_ (.A(_02424_),
    .B(_02427_),
    .Y(_02436_));
 sky130_fd_sc_hd__xor2_1 _08947_ (.A(_02435_),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _08948_ (.A0(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_02437_),
    .S(_02319_),
    .X(_02438_));
 sky130_fd_sc_hd__and2_1 _08949_ (.A(_01981_),
    .B(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__clkbuf_1 _08950_ (.A(_02439_),
    .X(_00274_));
 sky130_fd_sc_hd__a21boi_1 _08951_ (.A1(_02424_),
    .A2(_02427_),
    .B1_N(_02435_),
    .Y(_02440_));
 sky130_fd_sc_hd__inv_2 _08952_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_02441_));
 sky130_fd_sc_hd__or4_4 _08953_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .C(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .D(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__nand2_1 _08954_ (.A(_02342_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__xnor2_1 _08955_ (.A(_02441_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__and2_1 _08956_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__nor2_1 _08957_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_02444_),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_1 _08958_ (.A(_02445_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__o21a_1 _08959_ (.A1(_02433_),
    .A2(_02440_),
    .B1(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__nor3_1 _08960_ (.A(_02433_),
    .B(_02440_),
    .C(_02447_),
    .Y(_02449_));
 sky130_fd_sc_hd__o21ai_1 _08961_ (.A1(_02448_),
    .A2(_02449_),
    .B1(_02322_),
    .Y(_02450_));
 sky130_fd_sc_hd__o211a_1 _08962_ (.A1(_02321_),
    .A2(net486),
    .B1(_02381_),
    .C1(_02450_),
    .X(_00275_));
 sky130_fd_sc_hd__o21a_1 _08963_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A2(_02442_),
    .B1(_02341_),
    .X(_02451_));
 sky130_fd_sc_hd__xor2_2 _08964_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__xnor2_2 _08965_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__nor2_1 _08966_ (.A(_02445_),
    .B(_02448_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21oi_1 _08967_ (.A1(_02453_),
    .A2(_02454_),
    .B1(_02333_),
    .Y(_02455_));
 sky130_fd_sc_hd__o21ai_1 _08968_ (.A1(_02453_),
    .A2(_02454_),
    .B1(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__o211a_1 _08969_ (.A1(_02321_),
    .A2(net619),
    .B1(_02381_),
    .C1(_02456_),
    .X(_00276_));
 sky130_fd_sc_hd__and2_1 _08970_ (.A(_02448_),
    .B(_02453_),
    .X(_02457_));
 sky130_fd_sc_hd__inv_2 _08971_ (.A(_02452_),
    .Y(_02458_));
 sky130_fd_sc_hd__a21o_1 _08972_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_02458_),
    .B1(_02445_),
    .X(_02459_));
 sky130_fd_sc_hd__o21a_1 _08973_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_02458_),
    .B1(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__o31a_1 _08974_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A3(_02442_),
    .B1(_02342_),
    .X(_02461_));
 sky130_fd_sc_hd__xnor2_1 _08975_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_02461_),
    .Y(_02462_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__or2_1 _08977_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02462_),
    .X(_02464_));
 sky130_fd_sc_hd__and2_1 _08978_ (.A(_02463_),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__o21ai_1 _08979_ (.A1(_02457_),
    .A2(_02460_),
    .B1(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__o31a_1 _08980_ (.A1(_02465_),
    .A2(_02457_),
    .A3(_02460_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02467_));
 sky130_fd_sc_hd__a22o_1 _08981_ (.A1(_02313_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_02466_),
    .B2(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__and2_1 _08982_ (.A(_01981_),
    .B(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_1 _08983_ (.A(_02469_),
    .X(_00277_));
 sky130_fd_sc_hd__o41a_1 _08984_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A3(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A4(_02442_),
    .B1(_02341_),
    .X(_02470_));
 sky130_fd_sc_hd__xor2_1 _08985_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__or2b_1 _08986_ (.A(_02471_),
    .B_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_02472_));
 sky130_fd_sc_hd__inv_2 _08987_ (.A(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__and2b_1 _08988_ (.A_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_02471_),
    .X(_02474_));
 sky130_fd_sc_hd__nor2_1 _08989_ (.A(_02473_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__a21oi_1 _08990_ (.A1(_02463_),
    .A2(_02466_),
    .B1(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__a31o_1 _08991_ (.A1(_02463_),
    .A2(_02466_),
    .A3(_02475_),
    .B1(_02369_),
    .X(_02477_));
 sky130_fd_sc_hd__o221a_1 _08992_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_02476_),
    .B2(_02477_),
    .C1(_02414_),
    .X(_00278_));
 sky130_fd_sc_hd__o2111a_1 _08993_ (.A1(_02433_),
    .A2(_02440_),
    .B1(_02447_),
    .C1(_02453_),
    .D1(_02475_),
    .X(_02478_));
 sky130_fd_sc_hd__a21oi_1 _08994_ (.A1(_02463_),
    .A2(_02472_),
    .B1(_02474_),
    .Y(_02479_));
 sky130_fd_sc_hd__a31o_1 _08995_ (.A1(_02465_),
    .A2(_02460_),
    .A3(_02475_),
    .B1(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__a21o_1 _08996_ (.A1(_02465_),
    .A2(_02478_),
    .B1(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__or2_1 _08997_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_02482_));
 sky130_fd_sc_hd__or4_2 _08998_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .C(_02442_),
    .D(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__and2_1 _08999_ (.A(_02342_),
    .B(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__xnor2_1 _09000_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__or2_1 _09002_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02485_),
    .X(_02487_));
 sky130_fd_sc_hd__and2_1 _09003_ (.A(_02486_),
    .B(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__or2_1 _09004_ (.A(_02481_),
    .B(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(_02481_),
    .B(_02488_),
    .Y(_02490_));
 sky130_fd_sc_hd__a21o_1 _09006_ (.A1(_02489_),
    .A2(_02490_),
    .B1(_02333_),
    .X(_02491_));
 sky130_fd_sc_hd__o211a_1 _09007_ (.A1(_02321_),
    .A2(net616),
    .B1(_02381_),
    .C1(_02491_),
    .X(_00279_));
 sky130_fd_sc_hd__o21a_1 _09008_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_02483_),
    .B1(_02343_),
    .X(_02492_));
 sky130_fd_sc_hd__xor2_2 _09009_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__xnor2_1 _09010_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__a21oi_1 _09011_ (.A1(_02486_),
    .A2(_02490_),
    .B1(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__a31o_1 _09012_ (.A1(_02486_),
    .A2(_02490_),
    .A3(_02494_),
    .B1(_02369_),
    .X(_02496_));
 sky130_fd_sc_hd__o221a_1 _09013_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_02495_),
    .B2(_02496_),
    .C1(_02414_),
    .X(_00280_));
 sky130_fd_sc_hd__clkbuf_4 _09014_ (.A(_01765_),
    .X(_02497_));
 sky130_fd_sc_hd__inv_2 _09015_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .Y(_02498_));
 sky130_fd_sc_hd__o21a_1 _09016_ (.A1(_02498_),
    .A2(_02493_),
    .B1(_02486_),
    .X(_02499_));
 sky130_fd_sc_hd__a21o_1 _09017_ (.A1(_02498_),
    .A2(_02493_),
    .B1(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__nand2_1 _09018_ (.A(_02488_),
    .B(_02494_),
    .Y(_02501_));
 sky130_fd_sc_hd__inv_2 _09019_ (.A(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand2_1 _09020_ (.A(_02481_),
    .B(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__or3_1 _09021_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .C(_02483_),
    .X(_02504_));
 sky130_fd_sc_hd__and2_1 _09022_ (.A(_02343_),
    .B(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__xnor2_2 _09023_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__xor2_2 _09024_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__a21bo_1 _09025_ (.A1(_02500_),
    .A2(_02503_),
    .B1_N(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__nand3b_1 _09026_ (.A_N(_02507_),
    .B(_02500_),
    .C(_02503_),
    .Y(_02509_));
 sky130_fd_sc_hd__and2_1 _09027_ (.A(_02312_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_02510_));
 sky130_fd_sc_hd__a31o_1 _09028_ (.A1(_02319_),
    .A2(_02508_),
    .A3(_02509_),
    .B1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__and2_1 _09029_ (.A(_02497_),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _09030_ (.A(_02512_),
    .X(_00281_));
 sky130_fd_sc_hd__nand2_1 _09031_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02506_),
    .Y(_02513_));
 sky130_fd_sc_hd__o21a_1 _09032_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_02504_),
    .B1(_02343_),
    .X(_02514_));
 sky130_fd_sc_hd__xor2_2 _09033_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__xnor2_2 _09034_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__a21oi_1 _09035_ (.A1(_02513_),
    .A2(_02508_),
    .B1(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__a31o_1 _09036_ (.A1(_02513_),
    .A2(_02508_),
    .A3(_02516_),
    .B1(_02369_),
    .X(_02518_));
 sky130_fd_sc_hd__o221a_1 _09037_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_02517_),
    .B2(_02518_),
    .C1(_02414_),
    .X(_00282_));
 sky130_fd_sc_hd__and2_1 _09038_ (.A(_02507_),
    .B(_02516_),
    .X(_02519_));
 sky130_fd_sc_hd__inv_2 _09039_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .Y(_02520_));
 sky130_fd_sc_hd__nand2_1 _09040_ (.A(_02507_),
    .B(_02516_),
    .Y(_02521_));
 sky130_fd_sc_hd__a21o_1 _09041_ (.A1(_02520_),
    .A2(_02515_),
    .B1(_02513_),
    .X(_02522_));
 sky130_fd_sc_hd__o221ai_1 _09042_ (.A1(_02520_),
    .A2(_02515_),
    .B1(_02521_),
    .B2(_02500_),
    .C1(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__a31o_1 _09043_ (.A1(_02481_),
    .A2(_02502_),
    .A3(_02519_),
    .B1(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__or3_1 _09044_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .C(_02504_),
    .X(_02525_));
 sky130_fd_sc_hd__and2_1 _09045_ (.A(_02343_),
    .B(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__xnor2_1 _09046_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _09047_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__or2_1 _09048_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02527_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(_02528_),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__xnor2_1 _09050_ (.A(_02524_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__or2_1 _09051_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_02532_));
 sky130_fd_sc_hd__o211a_1 _09052_ (.A1(_02314_),
    .A2(_02531_),
    .B1(_02532_),
    .C1(_02260_),
    .X(_00283_));
 sky130_fd_sc_hd__or2b_1 _09053_ (.A(_02530_),
    .B_N(_02524_),
    .X(_02533_));
 sky130_fd_sc_hd__o21a_1 _09054_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_02525_),
    .B1(_02343_),
    .X(_02534_));
 sky130_fd_sc_hd__xor2_2 _09055_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__xnor2_1 _09056_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__a21oi_1 _09057_ (.A1(_02528_),
    .A2(_02533_),
    .B1(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__a31o_1 _09058_ (.A1(_02528_),
    .A2(_02533_),
    .A3(_02536_),
    .B1(_02369_),
    .X(_02538_));
 sky130_fd_sc_hd__o221a_1 _09059_ (.A1(_02387_),
    .A2(net644),
    .B1(_02537_),
    .B2(_02538_),
    .C1(_02414_),
    .X(_00284_));
 sky130_fd_sc_hd__or3_1 _09060_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .C(_02525_),
    .X(_02539_));
 sky130_fd_sc_hd__and2_1 _09061_ (.A(_02344_),
    .B(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__xnor2_1 _09062_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__xor2_1 _09063_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__and2b_1 _09064_ (.A_N(_02530_),
    .B(_02536_),
    .X(_02543_));
 sky130_fd_sc_hd__inv_2 _09065_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .Y(_02544_));
 sky130_fd_sc_hd__o21a_1 _09066_ (.A1(_02544_),
    .A2(_02535_),
    .B1(_02528_),
    .X(_02545_));
 sky130_fd_sc_hd__a21oi_1 _09067_ (.A1(_02544_),
    .A2(_02535_),
    .B1(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__a21o_1 _09068_ (.A1(_02524_),
    .A2(_02543_),
    .B1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_1 _09069_ (.A(_02542_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21a_1 _09070_ (.A1(_02542_),
    .A2(_02547_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02549_));
 sky130_fd_sc_hd__a22o_1 _09071_ (.A1(_02313_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_02548_),
    .B2(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__and2_1 _09072_ (.A(_02497_),
    .B(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_1 _09073_ (.A(_02551_),
    .X(_00285_));
 sky130_fd_sc_hd__nand2_1 _09074_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02541_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _09075_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02539_),
    .Y(_02553_));
 sky130_fd_sc_hd__or2_1 _09076_ (.A(_01958_),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_2 _09077_ (.A0(_02554_),
    .A1(_02344_),
    .S(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _09078_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_02553_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand3_1 _09079_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_02555_),
    .C(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__inv_2 _09080_ (.A(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__a21oi_1 _09081_ (.A1(_02555_),
    .A2(_02556_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _09082_ (.A(_02558_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__a21oi_1 _09083_ (.A1(_02552_),
    .A2(_02548_),
    .B1(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__a31o_1 _09084_ (.A1(_02552_),
    .A2(_02548_),
    .A3(_02560_),
    .B1(_02369_),
    .X(_02562_));
 sky130_fd_sc_hd__o221a_1 _09085_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B1(_02561_),
    .B2(_02562_),
    .C1(_02414_),
    .X(_00286_));
 sky130_fd_sc_hd__or2_1 _09086_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02555_),
    .X(_02563_));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02555_),
    .Y(_02564_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(_02563_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand2_1 _09089_ (.A(_02552_),
    .B(_02557_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_1 _09090_ (.A1(_02542_),
    .A2(_02547_),
    .B1(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__or3_1 _09091_ (.A(_02559_),
    .B(_02565_),
    .C(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__o21ai_1 _09092_ (.A1(_02559_),
    .A2(_02567_),
    .B1(_02565_),
    .Y(_02569_));
 sky130_fd_sc_hd__and2_1 _09093_ (.A(_02312_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .X(_02570_));
 sky130_fd_sc_hd__a31o_1 _09094_ (.A1(_02319_),
    .A2(_02568_),
    .A3(_02569_),
    .B1(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__and2_1 _09095_ (.A(_02497_),
    .B(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _09096_ (.A(_02572_),
    .X(_00287_));
 sky130_fd_sc_hd__xor2_1 _09097_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_02555_),
    .X(_02573_));
 sky130_fd_sc_hd__a21oi_1 _09098_ (.A1(_02564_),
    .A2(_02568_),
    .B1(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__a31o_1 _09099_ (.A1(_02564_),
    .A2(_02568_),
    .A3(_02573_),
    .B1(_02369_),
    .X(_02575_));
 sky130_fd_sc_hd__o221a_1 _09100_ (.A1(_02387_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B1(_02574_),
    .B2(_02575_),
    .C1(_02414_),
    .X(_00288_));
 sky130_fd_sc_hd__and2_1 _09101_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .X(_02576_));
 sky130_fd_sc_hd__nor2_1 _09102_ (.A(net273),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .Y(_02577_));
 sky130_fd_sc_hd__o21ai_1 _09103_ (.A1(_02576_),
    .A2(_02577_),
    .B1(_02322_),
    .Y(_02578_));
 sky130_fd_sc_hd__o211a_1 _09104_ (.A1(_02321_),
    .A2(net291),
    .B1(_02381_),
    .C1(_02578_),
    .X(_00289_));
 sky130_fd_sc_hd__and2b_1 _09105_ (.A_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .X(_02579_));
 sky130_fd_sc_hd__xnor2_1 _09106_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__xnor2_1 _09107_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__nor2_1 _09108_ (.A(_02576_),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__and2_1 _09109_ (.A(_02576_),
    .B(_02581_),
    .X(_02583_));
 sky130_fd_sc_hd__o21ai_1 _09110_ (.A1(_02582_),
    .A2(_02583_),
    .B1(_02320_),
    .Y(_02584_));
 sky130_fd_sc_hd__o211a_1 _09111_ (.A1(_02329_),
    .A2(net325),
    .B1(_02381_),
    .C1(_02584_),
    .X(_00290_));
 sky130_fd_sc_hd__and2b_1 _09112_ (.A_N(_02580_),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_02585_));
 sky130_fd_sc_hd__o21a_1 _09113_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_02341_),
    .X(_02586_));
 sky130_fd_sc_hd__xnor2_1 _09114_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__xnor2_1 _09115_ (.A(_02152_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__o21bai_2 _09116_ (.A1(_02585_),
    .A2(_02583_),
    .B1_N(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__or3b_1 _09117_ (.A(_02585_),
    .B(_02583_),
    .C_N(_02588_),
    .X(_02590_));
 sky130_fd_sc_hd__inv_2 _09118_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_02591_));
 sky130_fd_sc_hd__nor2_1 _09119_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__a31o_1 _09120_ (.A1(_02319_),
    .A2(_02589_),
    .A3(_02590_),
    .B1(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__and2_1 _09121_ (.A(_02497_),
    .B(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__clkbuf_1 _09122_ (.A(_02594_),
    .X(_00291_));
 sky130_fd_sc_hd__inv_2 _09123_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_02595_));
 sky130_fd_sc_hd__or2_1 _09124_ (.A(_02152_),
    .B(_02587_),
    .X(_02596_));
 sky130_fd_sc_hd__o31a_1 _09125_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A3(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_02341_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_1 _09126_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__nor2_1 _09127_ (.A(_02156_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__and2_1 _09128_ (.A(_02156_),
    .B(_02598_),
    .X(_02600_));
 sky130_fd_sc_hd__or2_1 _09129_ (.A(_02599_),
    .B(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__and3_1 _09130_ (.A(_02596_),
    .B(_02589_),
    .C(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__a21oi_2 _09131_ (.A1(_02596_),
    .A2(_02589_),
    .B1(_02601_),
    .Y(_02603_));
 sky130_fd_sc_hd__or3_1 _09132_ (.A(_02312_),
    .B(_02602_),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__o21a_1 _09133_ (.A1(_02319_),
    .A2(_02595_),
    .B1(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__and2b_1 _09134_ (.A_N(_02605_),
    .B(_01979_),
    .X(_02606_));
 sky130_fd_sc_hd__clkbuf_1 _09135_ (.A(_02606_),
    .X(_00292_));
 sky130_fd_sc_hd__inv_2 _09136_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_02607_));
 sky130_fd_sc_hd__or4_4 _09137_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .C(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .D(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .X(_02608_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(_02342_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__xor2_1 _09139_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__nor2_1 _09140_ (.A(_02607_),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__and2_1 _09141_ (.A(_02607_),
    .B(_02610_),
    .X(_02612_));
 sky130_fd_sc_hd__or2_1 _09142_ (.A(_02611_),
    .B(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__inv_2 _09143_ (.A(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__o21a_1 _09144_ (.A1(_02599_),
    .A2(_02603_),
    .B1(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__nor3_1 _09145_ (.A(_02599_),
    .B(_02603_),
    .C(_02614_),
    .Y(_02616_));
 sky130_fd_sc_hd__o21ai_1 _09146_ (.A1(_02615_),
    .A2(_02616_),
    .B1(_02320_),
    .Y(_02617_));
 sky130_fd_sc_hd__o211a_1 _09147_ (.A1(_02329_),
    .A2(net473),
    .B1(_02381_),
    .C1(_02617_),
    .X(_00293_));
 sky130_fd_sc_hd__o21a_1 _09148_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(_02608_),
    .B1(_02342_),
    .X(_02618_));
 sky130_fd_sc_hd__xor2_1 _09149_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__and2_1 _09150_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__or2_1 _09151_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_02619_),
    .X(_02621_));
 sky130_fd_sc_hd__and2b_1 _09152_ (.A_N(_02620_),
    .B(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__o21ba_1 _09153_ (.A1(_02611_),
    .A2(_02615_),
    .B1_N(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__or3b_1 _09154_ (.A(_02611_),
    .B(_02615_),
    .C_N(_02622_),
    .X(_02624_));
 sky130_fd_sc_hd__nand2_1 _09155_ (.A(_02320_),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__o221a_1 _09156_ (.A1(_02322_),
    .A2(net548),
    .B1(_02623_),
    .B2(_02625_),
    .C1(_02414_),
    .X(_00294_));
 sky130_fd_sc_hd__or2_1 _09157_ (.A(_02611_),
    .B(_02620_),
    .X(_02626_));
 sky130_fd_sc_hd__or2_1 _09158_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .X(_02627_));
 sky130_fd_sc_hd__o21a_1 _09159_ (.A1(_02608_),
    .A2(_02627_),
    .B1(_02342_),
    .X(_02628_));
 sky130_fd_sc_hd__xnor2_2 _09160_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__xnor2_2 _09161_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__o211ai_2 _09162_ (.A1(_02615_),
    .A2(_02626_),
    .B1(_02630_),
    .C1(_02621_),
    .Y(_02631_));
 sky130_fd_sc_hd__o211a_1 _09163_ (.A1(_02599_),
    .A2(_02603_),
    .B1(_02614_),
    .C1(_02622_),
    .X(_02632_));
 sky130_fd_sc_hd__a211o_1 _09164_ (.A1(_02621_),
    .A2(_02626_),
    .B1(_02632_),
    .C1(_02630_),
    .X(_02633_));
 sky130_fd_sc_hd__inv_2 _09165_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_02634_));
 sky130_fd_sc_hd__nor2_1 _09166_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__a31o_1 _09167_ (.A1(_02319_),
    .A2(_02631_),
    .A3(_02633_),
    .B1(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__and2_1 _09168_ (.A(_02497_),
    .B(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_1 _09169_ (.A(_02637_),
    .X(_00295_));
 sky130_fd_sc_hd__or2_1 _09170_ (.A(_02441_),
    .B(_02629_),
    .X(_02638_));
 sky130_fd_sc_hd__o31a_1 _09171_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_02608_),
    .A3(_02627_),
    .B1(_02342_),
    .X(_02639_));
 sky130_fd_sc_hd__xnor2_1 _09172_ (.A(_02498_),
    .B(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _09173_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__inv_2 _09174_ (.A(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__nor2_1 _09175_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02640_),
    .Y(_02643_));
 sky130_fd_sc_hd__nor2_1 _09176_ (.A(_02642_),
    .B(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__a21oi_1 _09177_ (.A1(_02638_),
    .A2(_02631_),
    .B1(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__a31o_1 _09178_ (.A1(_02638_),
    .A2(_02631_),
    .A3(_02644_),
    .B1(_02369_),
    .X(_02646_));
 sky130_fd_sc_hd__o221a_1 _09179_ (.A1(_02322_),
    .A2(net567),
    .B1(_02645_),
    .B2(_02646_),
    .C1(_02414_),
    .X(_00296_));
 sky130_fd_sc_hd__a21oi_1 _09180_ (.A1(_02638_),
    .A2(_02641_),
    .B1(_02643_),
    .Y(_02647_));
 sky130_fd_sc_hd__a41o_1 _09181_ (.A1(_02621_),
    .A2(_02630_),
    .A3(_02626_),
    .A4(_02644_),
    .B1(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__a31o_2 _09182_ (.A1(_02630_),
    .A2(_02632_),
    .A3(_02644_),
    .B1(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__inv_2 _09183_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_02650_));
 sky130_fd_sc_hd__or2_1 _09184_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_02651_));
 sky130_fd_sc_hd__or3_1 _09185_ (.A(_02608_),
    .B(_02627_),
    .C(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(_02342_),
    .B(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__xor2_1 _09187_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__nor2_1 _09188_ (.A(_02650_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__and2_1 _09189_ (.A(_02650_),
    .B(_02654_),
    .X(_02656_));
 sky130_fd_sc_hd__or2_1 _09190_ (.A(_02655_),
    .B(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__xnor2_1 _09191_ (.A(_02649_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__or2_1 _09192_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_02659_));
 sky130_fd_sc_hd__o211a_1 _09193_ (.A1(_02314_),
    .A2(_02658_),
    .B1(_02659_),
    .C1(_02260_),
    .X(_00297_));
 sky130_fd_sc_hd__o21a_1 _09194_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_02652_),
    .B1(_02342_),
    .X(_02660_));
 sky130_fd_sc_hd__xnor2_1 _09195_ (.A(_02520_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__and2_1 _09196_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__or2_1 _09197_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_02661_),
    .X(_02663_));
 sky130_fd_sc_hd__or2b_1 _09198_ (.A(_02662_),
    .B_N(_02663_),
    .X(_02664_));
 sky130_fd_sc_hd__and2b_1 _09199_ (.A_N(_02657_),
    .B(_02649_),
    .X(_02665_));
 sky130_fd_sc_hd__or2_1 _09200_ (.A(_02655_),
    .B(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__nor2_1 _09201_ (.A(_02664_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__a21o_1 _09202_ (.A1(_02664_),
    .A2(_02666_),
    .B1(_02333_),
    .X(_02668_));
 sky130_fd_sc_hd__o221a_1 _09203_ (.A1(_02322_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_02667_),
    .B2(_02668_),
    .C1(_02414_),
    .X(_00298_));
 sky130_fd_sc_hd__and2_1 _09204_ (.A(_02333_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .X(_02669_));
 sky130_fd_sc_hd__or2_1 _09205_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_02670_));
 sky130_fd_sc_hd__or4_1 _09206_ (.A(_02608_),
    .B(_02627_),
    .C(_02651_),
    .D(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__nand2_1 _09207_ (.A(_02343_),
    .B(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__xor2_1 _09208_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02672_),
    .X(_02673_));
 sky130_fd_sc_hd__or2_1 _09209_ (.A(_02237_),
    .B(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__nand2_1 _09210_ (.A(_02237_),
    .B(_02673_),
    .Y(_02675_));
 sky130_fd_sc_hd__nand2_1 _09211_ (.A(_02674_),
    .B(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__o21ai_1 _09212_ (.A1(_02655_),
    .A2(_02662_),
    .B1(_02663_),
    .Y(_02677_));
 sky130_fd_sc_hd__or2_1 _09213_ (.A(_02657_),
    .B(_02664_),
    .X(_02678_));
 sky130_fd_sc_hd__inv_2 _09214_ (.A(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_1 _09215_ (.A(_02649_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__a31o_1 _09216_ (.A1(_02676_),
    .A2(_02677_),
    .A3(_02680_),
    .B1(_02313_),
    .X(_02681_));
 sky130_fd_sc_hd__a21o_1 _09217_ (.A1(_02677_),
    .A2(_02680_),
    .B1(_02676_),
    .X(_02682_));
 sky130_fd_sc_hd__and2b_1 _09218_ (.A_N(_02681_),
    .B(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__o21a_1 _09219_ (.A1(_02669_),
    .A2(_02683_),
    .B1(_02132_),
    .X(_00299_));
 sky130_fd_sc_hd__o21a_1 _09220_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_02671_),
    .B1(_02343_),
    .X(_02684_));
 sky130_fd_sc_hd__xnor2_2 _09221_ (.A(_02544_),
    .B(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__xor2_1 _09222_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__a21oi_1 _09223_ (.A1(_02674_),
    .A2(_02682_),
    .B1(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__a31o_1 _09224_ (.A1(_02674_),
    .A2(_02682_),
    .A3(_02686_),
    .B1(_02313_),
    .X(_02688_));
 sky130_fd_sc_hd__buf_4 _09225_ (.A(_02308_),
    .X(_02689_));
 sky130_fd_sc_hd__o221a_1 _09226_ (.A1(_02322_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_02687_),
    .B2(_02688_),
    .C1(_02689_),
    .X(_00300_));
 sky130_fd_sc_hd__and2b_1 _09227_ (.A_N(_02676_),
    .B(_02686_),
    .X(_02690_));
 sky130_fd_sc_hd__o21a_1 _09228_ (.A1(_02655_),
    .A2(_02662_),
    .B1(_02663_),
    .X(_02691_));
 sky130_fd_sc_hd__o21ba_1 _09229_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_02685_),
    .B1_N(_02674_),
    .X(_02692_));
 sky130_fd_sc_hd__a221o_1 _09230_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_02685_),
    .B1(_02690_),
    .B2(_02691_),
    .C1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__a31o_1 _09231_ (.A1(_02649_),
    .A2(_02679_),
    .A3(_02690_),
    .B1(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__or3_1 _09232_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .C(_02671_),
    .X(_02695_));
 sky130_fd_sc_hd__and2_1 _09233_ (.A(_02343_),
    .B(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__xnor2_2 _09234_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__xor2_1 _09235_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__and2b_1 _09236_ (.A_N(_02694_),
    .B(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__and2b_1 _09237_ (.A_N(_02698_),
    .B(_02694_),
    .X(_02700_));
 sky130_fd_sc_hd__nor2_1 _09238_ (.A(_02699_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__or2_1 _09239_ (.A(_02315_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_02702_));
 sky130_fd_sc_hd__o211a_1 _09240_ (.A1(_02314_),
    .A2(_02701_),
    .B1(_02702_),
    .C1(_02260_),
    .X(_00301_));
 sky130_fd_sc_hd__o21a_1 _09241_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_02695_),
    .B1(_02343_),
    .X(_02703_));
 sky130_fd_sc_hd__xor2_2 _09242_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__xnor2_1 _09243_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__inv_2 _09244_ (.A(_02697_),
    .Y(_02706_));
 sky130_fd_sc_hd__a21o_1 _09245_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_02706_),
    .B1(_02700_),
    .X(_02707_));
 sky130_fd_sc_hd__o21ai_1 _09246_ (.A1(_02705_),
    .A2(_02707_),
    .B1(_02319_),
    .Y(_02708_));
 sky130_fd_sc_hd__a21o_1 _09247_ (.A1(_02705_),
    .A2(_02707_),
    .B1(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__o211a_1 _09248_ (.A1(_02329_),
    .A2(net534),
    .B1(_02381_),
    .C1(_02709_),
    .X(_00302_));
 sky130_fd_sc_hd__and2_1 _09249_ (.A(_02333_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_02710_));
 sky130_fd_sc_hd__inv_2 _09250_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .Y(_02711_));
 sky130_fd_sc_hd__nor3_1 _09251_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .C(_02695_),
    .Y(_02712_));
 sky130_fd_sc_hd__nor2_1 _09252_ (.A(_01958_),
    .B(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__xnor2_1 _09253_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__or2_1 _09254_ (.A(_02711_),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(_02711_),
    .B(_02714_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_1 _09256_ (.A(_02715_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__nor2_1 _09257_ (.A(_02698_),
    .B(_02705_),
    .Y(_02718_));
 sky130_fd_sc_hd__a22o_1 _09258_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_02706_),
    .B1(_02704_),
    .B2(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_02719_));
 sky130_fd_sc_hd__o21a_1 _09259_ (.A1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_02704_),
    .B1(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__a21oi_2 _09260_ (.A1(_02694_),
    .A2(_02718_),
    .B1(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__a21o_1 _09261_ (.A1(_02717_),
    .A2(_02721_),
    .B1(_02313_),
    .X(_02722_));
 sky130_fd_sc_hd__or2_1 _09262_ (.A(_02717_),
    .B(_02721_),
    .X(_02723_));
 sky130_fd_sc_hd__and2b_1 _09263_ (.A_N(_02722_),
    .B(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__o21a_1 _09264_ (.A1(_02710_),
    .A2(_02724_),
    .B1(_02132_),
    .X(_00303_));
 sky130_fd_sc_hd__a21oi_1 _09265_ (.A1(_02117_),
    .A2(_02712_),
    .B1(_01958_),
    .Y(_02725_));
 sky130_fd_sc_hd__mux2_2 _09266_ (.A0(_02725_),
    .A1(_01958_),
    .S(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_02726_));
 sky130_fd_sc_hd__and3_1 _09267_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_02117_),
    .C(_02712_),
    .X(_02727_));
 sky130_fd_sc_hd__o21ai_1 _09268_ (.A1(_02726_),
    .A2(_02727_),
    .B1(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .Y(_02728_));
 sky130_fd_sc_hd__or3_1 _09269_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_02726_),
    .C(_02727_),
    .X(_02729_));
 sky130_fd_sc_hd__nand2_1 _09270_ (.A(_02728_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__a21boi_1 _09271_ (.A1(_02715_),
    .A2(_02723_),
    .B1_N(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__a41o_1 _09272_ (.A1(_02715_),
    .A2(_02723_),
    .A3(_02728_),
    .A4(_02729_),
    .B1(_02313_),
    .X(_02732_));
 sky130_fd_sc_hd__o221a_1 _09273_ (.A1(_02322_),
    .A2(net579),
    .B1(_02731_),
    .B2(_02732_),
    .C1(_02689_),
    .X(_00304_));
 sky130_fd_sc_hd__xnor2_1 _09274_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02726_),
    .Y(_02733_));
 sky130_fd_sc_hd__a21bo_1 _09275_ (.A1(_02715_),
    .A2(_02728_),
    .B1_N(_02729_),
    .X(_02734_));
 sky130_fd_sc_hd__o31a_1 _09276_ (.A1(_02717_),
    .A2(_02721_),
    .A3(_02730_),
    .B1(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__nor2_1 _09277_ (.A(_02733_),
    .B(_02735_),
    .Y(_02736_));
 sky130_fd_sc_hd__a21o_1 _09278_ (.A1(_02733_),
    .A2(_02735_),
    .B1(_02312_),
    .X(_02737_));
 sky130_fd_sc_hd__o2bb2a_1 _09279_ (.A1_N(_02313_),
    .A2_N(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B1(_02736_),
    .B2(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__and2b_1 _09280_ (.A_N(_02738_),
    .B(_01979_),
    .X(_02739_));
 sky130_fd_sc_hd__clkbuf_1 _09281_ (.A(_02739_),
    .X(_00305_));
 sky130_fd_sc_hd__o2bb2a_1 _09282_ (.A1_N(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2_N(_02726_),
    .B1(_02733_),
    .B2(_02735_),
    .X(_02740_));
 sky130_fd_sc_hd__xnor2_1 _09283_ (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_02726_),
    .Y(_02741_));
 sky130_fd_sc_hd__xnor2_1 _09284_ (.A(_02740_),
    .B(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__o21ai_1 _09285_ (.A1(net626),
    .A2(_02320_),
    .B1(_01794_),
    .Y(_02743_));
 sky130_fd_sc_hd__a21oi_1 _09286_ (.A1(_02329_),
    .A2(_02742_),
    .B1(_02743_),
    .Y(_00306_));
 sky130_fd_sc_hd__and2_1 _09287_ (.A(_02320_),
    .B(_02310_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_1 _09288_ (.A(_02744_),
    .X(_00307_));
 sky130_fd_sc_hd__inv_2 _09289_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_02745_));
 sky130_fd_sc_hd__clkbuf_4 _09290_ (.A(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__buf_4 _09291_ (.A(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__clkbuf_4 _09292_ (.A(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__buf_4 _09293_ (.A(_01455_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_4 _09294_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02750_));
 sky130_fd_sc_hd__clkbuf_4 _09295_ (.A(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__or2_1 _09296_ (.A(net145),
    .B(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o211a_1 _09297_ (.A1(_02748_),
    .A2(net174),
    .B1(_02749_),
    .C1(_02752_),
    .X(_00308_));
 sky130_fd_sc_hd__or2_1 _09298_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_02751_),
    .X(_02753_));
 sky130_fd_sc_hd__o211a_1 _09299_ (.A1(_02748_),
    .A2(net210),
    .B1(_02749_),
    .C1(_02753_),
    .X(_00309_));
 sky130_fd_sc_hd__clkbuf_4 _09300_ (.A(_02751_),
    .X(_02754_));
 sky130_fd_sc_hd__clkbuf_4 _09301_ (.A(_02750_),
    .X(_02755_));
 sky130_fd_sc_hd__nand2_1 _09302_ (.A(_02755_),
    .B(net356),
    .Y(_02756_));
 sky130_fd_sc_hd__o211a_1 _09303_ (.A1(_02754_),
    .A2(net305),
    .B1(_02749_),
    .C1(_02756_),
    .X(_00310_));
 sky130_fd_sc_hd__clkbuf_4 _09304_ (.A(_02750_),
    .X(_02757_));
 sky130_fd_sc_hd__or2_1 _09305_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_02758_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .Y(_02759_));
 sky130_fd_sc_hd__a21oi_2 _09307_ (.A1(_02758_),
    .A2(_02759_),
    .B1(_02409_),
    .Y(_02760_));
 sky130_fd_sc_hd__buf_4 _09308_ (.A(_02746_),
    .X(_02761_));
 sky130_fd_sc_hd__a31o_1 _09309_ (.A1(_02409_),
    .A2(_02758_),
    .A3(_02759_),
    .B1(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__o221a_1 _09310_ (.A1(_02757_),
    .A2(net280),
    .B1(_02760_),
    .B2(_02762_),
    .C1(_02689_),
    .X(_00311_));
 sky130_fd_sc_hd__a21oi_1 _09311_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .Y(_02763_));
 sky130_fd_sc_hd__and3_1 _09312_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .C(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_02764_));
 sky130_fd_sc_hd__nor2_1 _09313_ (.A(_02763_),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_1 _09314_ (.A(_02760_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__a21o_1 _09315_ (.A1(_02760_),
    .A2(_02765_),
    .B1(_02747_),
    .X(_02767_));
 sky130_fd_sc_hd__o221a_1 _09316_ (.A1(_02757_),
    .A2(net313),
    .B1(_02766_),
    .B2(_02767_),
    .C1(_02689_),
    .X(_00312_));
 sky130_fd_sc_hd__and2_1 _09317_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(_02758_),
    .X(_02768_));
 sky130_fd_sc_hd__inv_2 _09318_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_02769_));
 sky130_fd_sc_hd__buf_2 _09319_ (.A(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__buf_2 _09320_ (.A(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__buf_4 _09321_ (.A(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _09322_ (.A0(_02763_),
    .A1(_02768_),
    .S(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__nor2_1 _09323_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__a21o_1 _09324_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(_02773_),
    .B1(_02747_),
    .X(_02775_));
 sky130_fd_sc_hd__o221a_1 _09325_ (.A1(_02757_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B1(_02774_),
    .B2(_02775_),
    .C1(_02689_),
    .X(_00313_));
 sky130_fd_sc_hd__a21o_1 _09326_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(_02776_));
 sky130_fd_sc_hd__or2_1 _09327_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_02768_),
    .X(_02777_));
 sky130_fd_sc_hd__nor2_1 _09328_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__a31o_1 _09329_ (.A1(_02409_),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A3(_02776_),
    .B1(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__and2_1 _09330_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__o21ai_1 _09331_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_02779_),
    .B1(_02755_),
    .Y(_02781_));
 sky130_fd_sc_hd__o221a_1 _09332_ (.A1(_02757_),
    .A2(net495),
    .B1(_02780_),
    .B2(_02781_),
    .C1(_02689_),
    .X(_00314_));
 sky130_fd_sc_hd__a21o_1 _09333_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_02777_),
    .B1(_02409_),
    .X(_02782_));
 sky130_fd_sc_hd__a21o_1 _09334_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(_02776_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(_02783_));
 sky130_fd_sc_hd__nand2_1 _09335_ (.A(_02409_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__inv_2 _09336_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .Y(_02785_));
 sky130_fd_sc_hd__a21oi_1 _09337_ (.A1(_02782_),
    .A2(_02784_),
    .B1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__a31o_1 _09338_ (.A1(_02785_),
    .A2(_02782_),
    .A3(_02784_),
    .B1(_02761_),
    .X(_02787_));
 sky130_fd_sc_hd__o221a_1 _09339_ (.A1(_02757_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B1(_02786_),
    .B2(_02787_),
    .C1(_02689_),
    .X(_00315_));
 sky130_fd_sc_hd__or2_1 _09340_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_02783_),
    .X(_02788_));
 sky130_fd_sc_hd__inv_2 _09341_ (.A(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__and3_1 _09342_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(_02777_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(_02789_),
    .A1(_02790_),
    .S(_02772_),
    .X(_02791_));
 sky130_fd_sc_hd__xnor2_1 _09344_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__nand2_1 _09345_ (.A(_02755_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__o211a_1 _09346_ (.A1(_02754_),
    .A2(net357),
    .B1(_02749_),
    .C1(_02793_),
    .X(_00316_));
 sky130_fd_sc_hd__or2_1 _09347_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_02788_),
    .X(_02794_));
 sky130_fd_sc_hd__inv_2 _09348_ (.A(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__and2_1 _09349_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_02790_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(_02795_),
    .A1(_02796_),
    .S(_02772_),
    .X(_02797_));
 sky130_fd_sc_hd__xnor2_1 _09351_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(_02755_),
    .B(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__o211a_1 _09353_ (.A1(_02754_),
    .A2(net395),
    .B1(_02749_),
    .C1(_02799_),
    .X(_00317_));
 sky130_fd_sc_hd__or2_1 _09354_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_02794_),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_1 _09355_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_02796_),
    .Y(_02801_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(_02800_),
    .A1(_02801_),
    .S(_02772_),
    .X(_02802_));
 sky130_fd_sc_hd__xnor2_1 _09357_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__buf_2 _09358_ (.A(_02750_),
    .X(_02804_));
 sky130_fd_sc_hd__or2_1 _09359_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(_02805_));
 sky130_fd_sc_hd__o211a_1 _09360_ (.A1(_02748_),
    .A2(_02803_),
    .B1(_02805_),
    .C1(_02260_),
    .X(_00318_));
 sky130_fd_sc_hd__and3_1 _09361_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .C(_02796_),
    .X(_02806_));
 sky130_fd_sc_hd__inv_2 _09362_ (.A(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__or2_1 _09363_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_02800_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(_02807_),
    .A1(_02808_),
    .S(_02409_),
    .X(_02809_));
 sky130_fd_sc_hd__and2_1 _09365_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__o21ai_1 _09366_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_02809_),
    .B1(_02755_),
    .Y(_02811_));
 sky130_fd_sc_hd__o221a_1 _09367_ (.A1(_02757_),
    .A2(net580),
    .B1(_02810_),
    .B2(_02811_),
    .C1(_02689_),
    .X(_00319_));
 sky130_fd_sc_hd__nand2_1 _09368_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_02806_),
    .Y(_02812_));
 sky130_fd_sc_hd__or2_1 _09369_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_02808_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(_02812_),
    .A1(_02813_),
    .S(_02409_),
    .X(_02814_));
 sky130_fd_sc_hd__and2_1 _09371_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__o21ai_1 _09372_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_02814_),
    .B1(_02751_),
    .Y(_02816_));
 sky130_fd_sc_hd__o221a_1 _09373_ (.A1(_02757_),
    .A2(net530),
    .B1(_02815_),
    .B2(_02816_),
    .C1(_02689_),
    .X(_00320_));
 sky130_fd_sc_hd__a31oi_2 _09374_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A3(_02806_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_02817_));
 sky130_fd_sc_hd__inv_2 _09375_ (.A(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__o21ai_1 _09376_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_02813_),
    .B1(_02409_),
    .Y(_02819_));
 sky130_fd_sc_hd__a21oi_1 _09377_ (.A1(_02818_),
    .A2(_02819_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .Y(_02820_));
 sky130_fd_sc_hd__a31o_1 _09378_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_02818_),
    .A3(_02819_),
    .B1(_02761_),
    .X(_02821_));
 sky130_fd_sc_hd__o221a_1 _09379_ (.A1(_02757_),
    .A2(net623),
    .B1(_02820_),
    .B2(_02821_),
    .C1(_02689_),
    .X(_00321_));
 sky130_fd_sc_hd__nand2_1 _09380_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_02819_),
    .Y(_02822_));
 sky130_fd_sc_hd__or2_1 _09381_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_02817_),
    .X(_02823_));
 sky130_fd_sc_hd__inv_2 _09382_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .Y(_02824_));
 sky130_fd_sc_hd__a21oi_1 _09383_ (.A1(_02822_),
    .A2(_02823_),
    .B1(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__a31o_1 _09384_ (.A1(_02824_),
    .A2(_02822_),
    .A3(_02823_),
    .B1(_02761_),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_4 _09385_ (.A(_02308_),
    .X(_02827_));
 sky130_fd_sc_hd__o221a_1 _09386_ (.A1(_02757_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_02825_),
    .B2(_02826_),
    .C1(_02827_),
    .X(_00322_));
 sky130_fd_sc_hd__inv_2 _09387_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .Y(_02828_));
 sky130_fd_sc_hd__o211a_1 _09388_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_02813_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(_02829_));
 sky130_fd_sc_hd__a311o_1 _09389_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A3(_02806_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(_02830_));
 sky130_fd_sc_hd__inv_2 _09390_ (.A(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(_02829_),
    .A1(_02831_),
    .S(_02772_),
    .X(_02832_));
 sky130_fd_sc_hd__a21oi_1 _09392_ (.A1(_02828_),
    .A2(_02832_),
    .B1(_02747_),
    .Y(_02833_));
 sky130_fd_sc_hd__o21ai_1 _09393_ (.A1(_02828_),
    .A2(_02832_),
    .B1(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__o211a_1 _09394_ (.A1(_02754_),
    .A2(net547),
    .B1(_02749_),
    .C1(_02834_),
    .X(_00323_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_02829_),
    .Y(_02835_));
 sky130_fd_sc_hd__or2_1 _09396_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_02830_),
    .X(_02836_));
 sky130_fd_sc_hd__mux2_1 _09397_ (.A0(_02835_),
    .A1(_02836_),
    .S(_02772_),
    .X(_02837_));
 sky130_fd_sc_hd__and2_1 _09398_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__o21ai_1 _09399_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_02837_),
    .B1(_02751_),
    .Y(_02839_));
 sky130_fd_sc_hd__o221a_1 _09400_ (.A1(_02757_),
    .A2(net601),
    .B1(_02838_),
    .B2(_02839_),
    .C1(_02827_),
    .X(_00324_));
 sky130_fd_sc_hd__xor2_1 _09401_ (.A(_02409_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(_02840_));
 sky130_fd_sc_hd__o21ai_1 _09402_ (.A1(_02837_),
    .A2(_02840_),
    .B1(net267),
    .Y(_02841_));
 sky130_fd_sc_hd__o31a_1 _09403_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_02837_),
    .A3(_02840_),
    .B1(_02751_),
    .X(_02842_));
 sky130_fd_sc_hd__o21ai_1 _09404_ (.A1(_02751_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_01794_),
    .Y(_02843_));
 sky130_fd_sc_hd__a21oi_1 _09405_ (.A1(_02841_),
    .A2(_02842_),
    .B1(_02843_),
    .Y(_00325_));
 sky130_fd_sc_hd__clkbuf_4 _09406_ (.A(_02750_),
    .X(_02844_));
 sky130_fd_sc_hd__o31ai_2 _09407_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_02836_),
    .B1(_02772_),
    .Y(_02845_));
 sky130_fd_sc_hd__a41o_1 _09408_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A4(_02829_),
    .B1(_02772_),
    .X(_02846_));
 sky130_fd_sc_hd__inv_2 _09409_ (.A(net440),
    .Y(_02847_));
 sky130_fd_sc_hd__a21oi_1 _09410_ (.A1(_02845_),
    .A2(_02846_),
    .B1(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__a31o_1 _09411_ (.A1(_02847_),
    .A2(_02845_),
    .A3(_02846_),
    .B1(_02761_),
    .X(_02849_));
 sky130_fd_sc_hd__o221a_1 _09412_ (.A1(_02844_),
    .A2(net474),
    .B1(_02848_),
    .B2(_02849_),
    .C1(_02827_),
    .X(_00326_));
 sky130_fd_sc_hd__buf_2 _09413_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_02850_));
 sky130_fd_sc_hd__buf_2 _09414_ (.A(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__nand2_1 _09415_ (.A(net440),
    .B(_02846_),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_1 _09416_ (.A1(_02845_),
    .A2(_02852_),
    .B1(_02747_),
    .X(_02853_));
 sky130_fd_sc_hd__o211a_1 _09417_ (.A1(_02754_),
    .A2(_02851_),
    .B1(_02749_),
    .C1(_02853_),
    .X(_00327_));
 sky130_fd_sc_hd__nor2_1 _09418_ (.A(_02595_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_02854_));
 sky130_fd_sc_hd__a21o_1 _09419_ (.A1(_02595_),
    .A2(net449),
    .B1(_02747_),
    .X(_02855_));
 sky130_fd_sc_hd__o221a_1 _09420_ (.A1(_02844_),
    .A2(net515),
    .B1(_02854_),
    .B2(_02855_),
    .C1(_02827_),
    .X(_00328_));
 sky130_fd_sc_hd__and2b_1 _09421_ (.A_N(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .X(_02856_));
 sky130_fd_sc_hd__xnor2_1 _09422_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__xnor2_1 _09423_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__xor2_1 _09424_ (.A(_02854_),
    .B(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__or2_1 _09425_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_02860_));
 sky130_fd_sc_hd__o211a_1 _09426_ (.A1(_02748_),
    .A2(_02859_),
    .B1(_02860_),
    .C1(_02260_),
    .X(_00329_));
 sky130_fd_sc_hd__and2_1 _09427_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_02857_),
    .X(_02861_));
 sky130_fd_sc_hd__nor2_1 _09428_ (.A(_02854_),
    .B(_02858_),
    .Y(_02862_));
 sky130_fd_sc_hd__o21ba_1 _09429_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B1_N(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_02863_));
 sky130_fd_sc_hd__xnor2_1 _09430_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__or2_1 _09431_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_02864_),
    .Y(_02866_));
 sky130_fd_sc_hd__and2_1 _09433_ (.A(_02865_),
    .B(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__o21ai_2 _09434_ (.A1(_02861_),
    .A2(_02862_),
    .B1(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__o31a_1 _09435_ (.A1(_02861_),
    .A2(_02862_),
    .A3(_02867_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02869_));
 sky130_fd_sc_hd__a22oi_1 _09436_ (.A1(_02746_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_02868_),
    .B2(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__and2b_1 _09437_ (.A_N(_02870_),
    .B(_01979_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_1 _09438_ (.A(_02871_),
    .X(_00330_));
 sky130_fd_sc_hd__o31a_1 _09439_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A3(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B1(_02769_),
    .X(_02872_));
 sky130_fd_sc_hd__xnor2_1 _09440_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__and2_1 _09441_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__nor2_1 _09442_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_02873_),
    .Y(_02875_));
 sky130_fd_sc_hd__nor2_1 _09443_ (.A(_02874_),
    .B(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_02866_),
    .B(_02868_),
    .Y(_02877_));
 sky130_fd_sc_hd__xor2_1 _09445_ (.A(_02876_),
    .B(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _09446_ (.A0(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_02878_),
    .S(_02750_),
    .X(_02879_));
 sky130_fd_sc_hd__and2_1 _09447_ (.A(_02497_),
    .B(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__clkbuf_1 _09448_ (.A(_02880_),
    .X(_00331_));
 sky130_fd_sc_hd__a21boi_1 _09449_ (.A1(_02866_),
    .A2(_02868_),
    .B1_N(_02876_),
    .Y(_02881_));
 sky130_fd_sc_hd__or4_2 _09450_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .C(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .D(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .X(_02882_));
 sky130_fd_sc_hd__nand2_1 _09451_ (.A(_02770_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__xor2_1 _09452_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__and2_1 _09453_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__nor2_1 _09454_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_02884_),
    .Y(_02886_));
 sky130_fd_sc_hd__nor2_1 _09455_ (.A(_02885_),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__o21a_1 _09456_ (.A1(_02874_),
    .A2(_02881_),
    .B1(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__nor3_1 _09457_ (.A(_02874_),
    .B(_02881_),
    .C(_02887_),
    .Y(_02889_));
 sky130_fd_sc_hd__o21ai_1 _09458_ (.A1(_02888_),
    .A2(_02889_),
    .B1(_02755_),
    .Y(_02890_));
 sky130_fd_sc_hd__o211a_1 _09459_ (.A1(_02754_),
    .A2(net527),
    .B1(_02749_),
    .C1(_02890_),
    .X(_00332_));
 sky130_fd_sc_hd__inv_2 _09460_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_02891_));
 sky130_fd_sc_hd__o21a_1 _09461_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(_02882_),
    .B1(_02769_),
    .X(_02892_));
 sky130_fd_sc_hd__xnor2_2 _09462_ (.A(_02891_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__xor2_2 _09463_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__o21a_1 _09464_ (.A1(_02885_),
    .A2(_02888_),
    .B1(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__o31ai_1 _09465_ (.A1(_02885_),
    .A2(_02888_),
    .A3(_02894_),
    .B1(_02751_),
    .Y(_02896_));
 sky130_fd_sc_hd__o221a_1 _09466_ (.A1(_02844_),
    .A2(net585),
    .B1(_02895_),
    .B2(_02896_),
    .C1(_02827_),
    .X(_00333_));
 sky130_fd_sc_hd__inv_2 _09467_ (.A(_02894_),
    .Y(_02897_));
 sky130_fd_sc_hd__and2_1 _09468_ (.A(_02888_),
    .B(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__inv_2 _09469_ (.A(_02893_),
    .Y(_02899_));
 sky130_fd_sc_hd__a21o_1 _09470_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_02899_),
    .B1(_02885_),
    .X(_02900_));
 sky130_fd_sc_hd__o21a_1 _09471_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_02899_),
    .B1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__or3_1 _09472_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .C(_02882_),
    .X(_02902_));
 sky130_fd_sc_hd__and2_1 _09473_ (.A(_02770_),
    .B(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__xnor2_1 _09474_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_1 _09475_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__or2_1 _09476_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_02904_),
    .X(_02906_));
 sky130_fd_sc_hd__and2_1 _09477_ (.A(_02905_),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__o21ai_1 _09478_ (.A1(_02898_),
    .A2(_02901_),
    .B1(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__o31a_1 _09479_ (.A1(_02907_),
    .A2(_02898_),
    .A3(_02901_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02909_));
 sky130_fd_sc_hd__a22o_1 _09480_ (.A1(_02746_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_02908_),
    .B2(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__and2_1 _09481_ (.A(_02497_),
    .B(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _09482_ (.A(_02911_),
    .X(_00334_));
 sky130_fd_sc_hd__o21a_1 _09483_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_02902_),
    .B1(_02770_),
    .X(_02912_));
 sky130_fd_sc_hd__xor2_2 _09484_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__xnor2_2 _09485_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__a21oi_1 _09486_ (.A1(_02905_),
    .A2(_02908_),
    .B1(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__a31o_1 _09487_ (.A1(_02905_),
    .A2(_02908_),
    .A3(_02914_),
    .B1(_02761_),
    .X(_02916_));
 sky130_fd_sc_hd__o221a_1 _09488_ (.A1(_02844_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_02915_),
    .B2(_02916_),
    .C1(_02827_),
    .X(_00335_));
 sky130_fd_sc_hd__or2_1 _09489_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_02917_));
 sky130_fd_sc_hd__or4_2 _09490_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .C(_02882_),
    .D(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__nand2_1 _09491_ (.A(_02771_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__xor2_1 _09492_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__nand2_1 _09493_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__or2_1 _09494_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_02920_),
    .X(_02922_));
 sky130_fd_sc_hd__and2_1 _09495_ (.A(_02921_),
    .B(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__inv_2 _09496_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .Y(_02924_));
 sky130_fd_sc_hd__o21ai_1 _09497_ (.A1(_02924_),
    .A2(_02913_),
    .B1(_02905_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _09498_ (.A(_02924_),
    .B(_02913_),
    .Y(_02926_));
 sky130_fd_sc_hd__a32o_1 _09499_ (.A1(_02907_),
    .A2(_02901_),
    .A3(_02914_),
    .B1(_02925_),
    .B2(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__a31o_1 _09500_ (.A1(_02907_),
    .A2(_02898_),
    .A3(_02914_),
    .B1(_02927_),
    .X(_02928_));
 sky130_fd_sc_hd__or2_1 _09501_ (.A(_02923_),
    .B(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__nand2_1 _09502_ (.A(_02923_),
    .B(_02928_),
    .Y(_02930_));
 sky130_fd_sc_hd__a21o_1 _09503_ (.A1(_02929_),
    .A2(_02930_),
    .B1(_02747_),
    .X(_02931_));
 sky130_fd_sc_hd__o211a_1 _09504_ (.A1(_02754_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_02749_),
    .C1(_02931_),
    .X(_00336_));
 sky130_fd_sc_hd__o21a_1 _09505_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_02918_),
    .B1(_02771_),
    .X(_02932_));
 sky130_fd_sc_hd__xor2_2 _09506_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__xnor2_1 _09507_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__a21oi_1 _09508_ (.A1(_02921_),
    .A2(_02930_),
    .B1(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__a31o_1 _09509_ (.A1(_02921_),
    .A2(_02930_),
    .A3(_02934_),
    .B1(_02761_),
    .X(_02936_));
 sky130_fd_sc_hd__o221a_1 _09510_ (.A1(_02844_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_02935_),
    .B2(_02936_),
    .C1(_02827_),
    .X(_00337_));
 sky130_fd_sc_hd__o31a_1 _09511_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A3(_02918_),
    .B1(_02771_),
    .X(_02937_));
 sky130_fd_sc_hd__xnor2_1 _09512_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__xor2_1 _09513_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(_02923_),
    .B(_02934_),
    .Y(_02940_));
 sky130_fd_sc_hd__inv_2 _09515_ (.A(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__inv_2 _09516_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .Y(_02942_));
 sky130_fd_sc_hd__o21a_1 _09517_ (.A1(_02942_),
    .A2(_02933_),
    .B1(_02921_),
    .X(_02943_));
 sky130_fd_sc_hd__a21o_1 _09518_ (.A1(_02942_),
    .A2(_02933_),
    .B1(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__a21bo_1 _09519_ (.A1(_02928_),
    .A2(_02941_),
    .B1_N(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(_02939_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__o21a_1 _09521_ (.A1(_02939_),
    .A2(_02945_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_02947_));
 sky130_fd_sc_hd__a22o_1 _09522_ (.A1(_02746_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_02946_),
    .B2(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__and2_1 _09523_ (.A(_02497_),
    .B(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _09524_ (.A(_02949_),
    .X(_00338_));
 sky130_fd_sc_hd__nand2_1 _09525_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_02938_),
    .Y(_02950_));
 sky130_fd_sc_hd__a21o_1 _09526_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_02771_),
    .B1(_02937_),
    .X(_02951_));
 sky130_fd_sc_hd__xor2_2 _09527_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__xnor2_1 _09528_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__a21oi_1 _09529_ (.A1(_02950_),
    .A2(_02946_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__a31o_1 _09530_ (.A1(_02950_),
    .A2(_02946_),
    .A3(_02953_),
    .B1(_02761_),
    .X(_02955_));
 sky130_fd_sc_hd__o221a_1 _09531_ (.A1(_02844_),
    .A2(net521),
    .B1(_02954_),
    .B2(_02955_),
    .C1(_02827_),
    .X(_00339_));
 sky130_fd_sc_hd__inv_2 _09532_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .Y(_02956_));
 sky130_fd_sc_hd__nand2_1 _09533_ (.A(_02956_),
    .B(_02952_),
    .Y(_02957_));
 sky130_fd_sc_hd__o21ai_1 _09534_ (.A1(_02956_),
    .A2(_02952_),
    .B1(_02950_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_02939_),
    .B(_02953_),
    .Y(_02959_));
 sky130_fd_sc_hd__nor2_1 _09536_ (.A(_02940_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__nor2_1 _09537_ (.A(_02944_),
    .B(_02959_),
    .Y(_02961_));
 sky130_fd_sc_hd__a221o_2 _09538_ (.A1(_02957_),
    .A2(_02958_),
    .B1(_02960_),
    .B2(_02928_),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__or2_1 _09539_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_02963_));
 sky130_fd_sc_hd__or4_4 _09540_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .C(_02918_),
    .D(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__and2_1 _09541_ (.A(_02771_),
    .B(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__xnor2_1 _09542_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__or2_1 _09544_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_02966_),
    .X(_02968_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_02967_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__xnor2_1 _09546_ (.A(_02962_),
    .B(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__or2_1 _09547_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_02971_));
 sky130_fd_sc_hd__o211a_1 _09548_ (.A1(_02748_),
    .A2(_02970_),
    .B1(_02971_),
    .C1(_02260_),
    .X(_00340_));
 sky130_fd_sc_hd__inv_2 _09549_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .Y(_02972_));
 sky130_fd_sc_hd__o21a_1 _09550_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(_02964_),
    .B1(_02772_),
    .X(_02973_));
 sky130_fd_sc_hd__xor2_2 _09551_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__xnor2_1 _09552_ (.A(_02972_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__inv_2 _09553_ (.A(_02969_),
    .Y(_02976_));
 sky130_fd_sc_hd__a21bo_1 _09554_ (.A1(_02962_),
    .A2(_02976_),
    .B1_N(_02967_),
    .X(_02977_));
 sky130_fd_sc_hd__nor2_1 _09555_ (.A(_02975_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__a21o_1 _09556_ (.A1(_02975_),
    .A2(_02977_),
    .B1(_02747_),
    .X(_02979_));
 sky130_fd_sc_hd__o221a_1 _09557_ (.A1(_02844_),
    .A2(net636),
    .B1(_02978_),
    .B2(_02979_),
    .C1(_02827_),
    .X(_00341_));
 sky130_fd_sc_hd__o21a_1 _09558_ (.A1(_02972_),
    .A2(_02974_),
    .B1(_02967_),
    .X(_02980_));
 sky130_fd_sc_hd__a21o_1 _09559_ (.A1(_02972_),
    .A2(_02974_),
    .B1(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__nor2_1 _09560_ (.A(_02969_),
    .B(_02975_),
    .Y(_02982_));
 sky130_fd_sc_hd__nand2_1 _09561_ (.A(_02962_),
    .B(_02982_),
    .Y(_02983_));
 sky130_fd_sc_hd__nor3_2 _09562_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .C(_02964_),
    .Y(_02984_));
 sky130_fd_sc_hd__or2_1 _09563_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_2 _09564_ (.A0(_02985_),
    .A1(_02771_),
    .S(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_02986_));
 sky130_fd_sc_hd__a21boi_2 _09565_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_02984_),
    .B1_N(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__xnor2_2 _09566_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__a21o_1 _09567_ (.A1(_02981_),
    .A2(_02983_),
    .B1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__a31oi_1 _09568_ (.A1(_02988_),
    .A2(_02981_),
    .A3(_02983_),
    .B1(_02745_),
    .Y(_02990_));
 sky130_fd_sc_hd__a22o_1 _09569_ (.A1(_02746_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_02989_),
    .B2(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__and2_1 _09570_ (.A(_02497_),
    .B(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _09571_ (.A(_02992_),
    .X(_00342_));
 sky130_fd_sc_hd__nand2_1 _09572_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_02987_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand2_1 _09573_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_02986_),
    .Y(_02994_));
 sky130_fd_sc_hd__or2_1 _09574_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_02986_),
    .X(_02995_));
 sky130_fd_sc_hd__and2_1 _09575_ (.A(_02994_),
    .B(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__a21oi_1 _09576_ (.A1(_02993_),
    .A2(_02989_),
    .B1(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__a31o_1 _09577_ (.A1(_02993_),
    .A2(_02989_),
    .A3(_02996_),
    .B1(_02761_),
    .X(_02998_));
 sky130_fd_sc_hd__o221a_1 _09578_ (.A1(_02844_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B1(_02997_),
    .B2(_02998_),
    .C1(_02827_),
    .X(_00343_));
 sky130_fd_sc_hd__or2_1 _09579_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02986_),
    .X(_02999_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_02986_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2_1 _09581_ (.A(_02999_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__and3b_1 _09582_ (.A_N(_02988_),
    .B(_02982_),
    .C(_02996_),
    .X(_03002_));
 sky130_fd_sc_hd__or2b_1 _09583_ (.A(_02988_),
    .B_N(_02996_),
    .X(_03003_));
 sky130_fd_sc_hd__o211a_1 _09584_ (.A1(_02981_),
    .A2(_03003_),
    .B1(_02994_),
    .C1(_02993_),
    .X(_03004_));
 sky130_fd_sc_hd__a21bo_1 _09585_ (.A1(_02962_),
    .A2(_03002_),
    .B1_N(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__xnor2_1 _09586_ (.A(_03001_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A1(_03006_),
    .S(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03007_));
 sky130_fd_sc_hd__and2_1 _09588_ (.A(_02497_),
    .B(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _09589_ (.A(_03008_),
    .X(_00344_));
 sky130_fd_sc_hd__or2b_1 _09590_ (.A(_03001_),
    .B_N(_03005_),
    .X(_03009_));
 sky130_fd_sc_hd__xor2_1 _09591_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_02986_),
    .X(_03010_));
 sky130_fd_sc_hd__a21oi_1 _09592_ (.A1(_03000_),
    .A2(_03009_),
    .B1(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__a31o_1 _09593_ (.A1(_03000_),
    .A2(_03009_),
    .A3(_03010_),
    .B1(_02746_),
    .X(_03012_));
 sky130_fd_sc_hd__buf_4 _09594_ (.A(_02308_),
    .X(_03013_));
 sky130_fd_sc_hd__o221a_1 _09595_ (.A1(_02844_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B1(_03011_),
    .B2(_03012_),
    .C1(_03013_),
    .X(_00345_));
 sky130_fd_sc_hd__and2_1 _09596_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .X(_03014_));
 sky130_fd_sc_hd__nor2_1 _09597_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .Y(_03015_));
 sky130_fd_sc_hd__o21ai_1 _09598_ (.A1(_03014_),
    .A2(_03015_),
    .B1(_02755_),
    .Y(_03016_));
 sky130_fd_sc_hd__o211a_1 _09599_ (.A1(_02754_),
    .A2(net478),
    .B1(_02749_),
    .C1(_03016_),
    .X(_00346_));
 sky130_fd_sc_hd__buf_4 _09600_ (.A(_01455_),
    .X(_03017_));
 sky130_fd_sc_hd__and2b_1 _09601_ (.A_N(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .X(_03018_));
 sky130_fd_sc_hd__xnor2_1 _09602_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__xnor2_1 _09603_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__nor2_1 _09604_ (.A(_03014_),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__and2_1 _09605_ (.A(_03014_),
    .B(_03020_),
    .X(_03022_));
 sky130_fd_sc_hd__o21ai_1 _09606_ (.A1(_03021_),
    .A2(_03022_),
    .B1(_02755_),
    .Y(_03023_));
 sky130_fd_sc_hd__o211a_1 _09607_ (.A1(_02754_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B1(_03017_),
    .C1(_03023_),
    .X(_00347_));
 sky130_fd_sc_hd__clkbuf_4 _09608_ (.A(_01765_),
    .X(_03024_));
 sky130_fd_sc_hd__and2b_1 _09609_ (.A_N(_03019_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_03025_));
 sky130_fd_sc_hd__o21a_1 _09610_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B1(_02769_),
    .X(_03026_));
 sky130_fd_sc_hd__xnor2_1 _09611_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__xnor2_1 _09612_ (.A(_02591_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__o21bai_2 _09613_ (.A1(_03025_),
    .A2(_03022_),
    .B1_N(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__or3b_1 _09614_ (.A(_03025_),
    .B(_03022_),
    .C_N(_03028_),
    .X(_03030_));
 sky130_fd_sc_hd__inv_2 _09615_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2_1 _09616_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__a31o_1 _09617_ (.A1(_02750_),
    .A2(_03029_),
    .A3(_03030_),
    .B1(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__and2_1 _09618_ (.A(_03024_),
    .B(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _09619_ (.A(_03034_),
    .X(_00348_));
 sky130_fd_sc_hd__inv_2 _09620_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_03035_));
 sky130_fd_sc_hd__or2_1 _09621_ (.A(_02591_),
    .B(_03027_),
    .X(_03036_));
 sky130_fd_sc_hd__o31a_1 _09622_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A3(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B1(_02769_),
    .X(_03037_));
 sky130_fd_sc_hd__xnor2_1 _09623_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__nor2_1 _09624_ (.A(_02595_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__and2_1 _09625_ (.A(_02595_),
    .B(_03038_),
    .X(_03040_));
 sky130_fd_sc_hd__or2_1 _09626_ (.A(_03039_),
    .B(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__and3_1 _09627_ (.A(_03036_),
    .B(_03029_),
    .C(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__a21oi_2 _09628_ (.A1(_03036_),
    .A2(_03029_),
    .B1(_03041_),
    .Y(_03043_));
 sky130_fd_sc_hd__or3_1 _09629_ (.A(_02745_),
    .B(_03042_),
    .C(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__o21a_1 _09630_ (.A1(_02750_),
    .A2(_03035_),
    .B1(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__and2b_1 _09631_ (.A_N(_03045_),
    .B(_01979_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _09632_ (.A(_03046_),
    .X(_00349_));
 sky130_fd_sc_hd__inv_2 _09633_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_03047_));
 sky130_fd_sc_hd__or4_2 _09634_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .C(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .D(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .X(_03048_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_02770_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__xnor2_1 _09636_ (.A(_02924_),
    .B(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2_1 _09637_ (.A(_03047_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__and2_1 _09638_ (.A(_03047_),
    .B(_03050_),
    .X(_03052_));
 sky130_fd_sc_hd__nor2_1 _09639_ (.A(_03051_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__o21a_1 _09640_ (.A1(_03039_),
    .A2(_03043_),
    .B1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__nor3_1 _09641_ (.A(_03039_),
    .B(_03043_),
    .C(_03053_),
    .Y(_03055_));
 sky130_fd_sc_hd__nor2_1 _09642_ (.A(_03054_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__or2_1 _09643_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_03057_));
 sky130_fd_sc_hd__buf_4 _09644_ (.A(_01474_),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _09645_ (.A1(_02748_),
    .A2(_03056_),
    .B1(_03057_),
    .C1(_03058_),
    .X(_00350_));
 sky130_fd_sc_hd__o21a_1 _09646_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(_03048_),
    .B1(_02770_),
    .X(_03059_));
 sky130_fd_sc_hd__xor2_1 _09647_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__and2_1 _09648_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__nor2_1 _09649_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03060_),
    .Y(_03062_));
 sky130_fd_sc_hd__nor2_2 _09650_ (.A(_03061_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__nor2_1 _09651_ (.A(_03051_),
    .B(_03054_),
    .Y(_03064_));
 sky130_fd_sc_hd__nor2_1 _09652_ (.A(_03063_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__a21o_1 _09653_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_02747_),
    .X(_03066_));
 sky130_fd_sc_hd__o221a_1 _09654_ (.A1(_02844_),
    .A2(net573),
    .B1(_03065_),
    .B2(_03066_),
    .C1(_03013_),
    .X(_00351_));
 sky130_fd_sc_hd__nor2_1 _09655_ (.A(_03062_),
    .B(_03064_),
    .Y(_03067_));
 sky130_fd_sc_hd__or2_1 _09656_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_03068_));
 sky130_fd_sc_hd__or2_1 _09657_ (.A(_03048_),
    .B(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__and2_1 _09658_ (.A(_02770_),
    .B(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__xnor2_1 _09659_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__or2_1 _09660_ (.A(_02634_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__nand2_1 _09661_ (.A(_02634_),
    .B(_03071_),
    .Y(_03073_));
 sky130_fd_sc_hd__and2_2 _09662_ (.A(_03072_),
    .B(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__o21ai_2 _09663_ (.A1(_03061_),
    .A2(_03067_),
    .B1(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__o31a_1 _09664_ (.A1(_03061_),
    .A2(_03067_),
    .A3(_03074_),
    .B1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03076_));
 sky130_fd_sc_hd__a22o_1 _09665_ (.A1(_02746_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1(_03075_),
    .B2(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__and2_1 _09666_ (.A(_03024_),
    .B(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _09667_ (.A(_03078_),
    .X(_00352_));
 sky130_fd_sc_hd__o21a_1 _09668_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_03069_),
    .B1(_02770_),
    .X(_03079_));
 sky130_fd_sc_hd__xor2_1 _09669_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__or2_1 _09671_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03080_),
    .X(_03082_));
 sky130_fd_sc_hd__and2_2 _09672_ (.A(_03081_),
    .B(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__a21oi_1 _09673_ (.A1(_03072_),
    .A2(_03075_),
    .B1(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__a31o_1 _09674_ (.A1(_03072_),
    .A2(_03075_),
    .A3(_03083_),
    .B1(_02746_),
    .X(_03085_));
 sky130_fd_sc_hd__o221a_1 _09675_ (.A1(_02755_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B1(_03084_),
    .B2(_03085_),
    .C1(_03013_),
    .X(_00353_));
 sky130_fd_sc_hd__or2_1 _09676_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_03086_));
 sky130_fd_sc_hd__or2_1 _09677_ (.A(_03069_),
    .B(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__nand2_1 _09678_ (.A(_02771_),
    .B(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__xor2_1 _09679_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__xnor2_1 _09680_ (.A(_02891_),
    .B(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__o21ba_1 _09681_ (.A1(_03051_),
    .A2(_03061_),
    .B1_N(_03062_),
    .X(_03091_));
 sky130_fd_sc_hd__nand2_1 _09682_ (.A(_03072_),
    .B(_03081_),
    .Y(_03092_));
 sky130_fd_sc_hd__a32o_1 _09683_ (.A1(_03074_),
    .A2(_03091_),
    .A3(_03083_),
    .B1(_03092_),
    .B2(_03082_),
    .X(_03093_));
 sky130_fd_sc_hd__a41o_1 _09684_ (.A1(_03054_),
    .A2(_03063_),
    .A3(_03074_),
    .A4(_03083_),
    .B1(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__xnor2_1 _09685_ (.A(_03090_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__or2_1 _09686_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_03096_));
 sky130_fd_sc_hd__o211a_1 _09687_ (.A1(_02748_),
    .A2(_03095_),
    .B1(_03096_),
    .C1(_03058_),
    .X(_00354_));
 sky130_fd_sc_hd__o21a_1 _09688_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_03087_),
    .B1(_02770_),
    .X(_03097_));
 sky130_fd_sc_hd__xor2_2 _09689_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__xnor2_1 _09690_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__a41oi_4 _09691_ (.A1(_03054_),
    .A2(_03063_),
    .A3(_03074_),
    .A4(_03083_),
    .B1(_03093_),
    .Y(_03100_));
 sky130_fd_sc_hd__or2_1 _09692_ (.A(_02891_),
    .B(_03089_),
    .X(_03101_));
 sky130_fd_sc_hd__o21ai_1 _09693_ (.A1(_03090_),
    .A2(_03100_),
    .B1(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__xnor2_1 _09694_ (.A(_03099_),
    .B(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__or2_1 _09695_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_03104_));
 sky130_fd_sc_hd__o211a_1 _09696_ (.A1(_02748_),
    .A2(_03103_),
    .B1(_03104_),
    .C1(_03058_),
    .X(_00355_));
 sky130_fd_sc_hd__inv_2 _09697_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .Y(_03105_));
 sky130_fd_sc_hd__or2_1 _09698_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_03106_));
 sky130_fd_sc_hd__or4_1 _09699_ (.A(_03048_),
    .B(_03068_),
    .C(_03086_),
    .D(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__nand2_1 _09700_ (.A(_02771_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__xnor2_2 _09701_ (.A(_02972_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__xor2_2 _09702_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__or2_1 _09703_ (.A(_03090_),
    .B(_03099_),
    .X(_03111_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03098_),
    .Y(_03112_));
 sky130_fd_sc_hd__nor2_1 _09705_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03098_),
    .Y(_03113_));
 sky130_fd_sc_hd__a21o_1 _09706_ (.A1(_03101_),
    .A2(_03112_),
    .B1(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__o21a_1 _09707_ (.A1(_03100_),
    .A2(_03111_),
    .B1(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__xnor2_1 _09708_ (.A(_03110_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__mux2_1 _09709_ (.A0(_03105_),
    .A1(_03116_),
    .S(_02750_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_6 _09710_ (.A(_01765_),
    .X(_03118_));
 sky130_fd_sc_hd__and2b_1 _09711_ (.A_N(_03117_),
    .B(_03118_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _09712_ (.A(_03119_),
    .X(_00356_));
 sky130_fd_sc_hd__o21a_1 _09713_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_03107_),
    .B1(_02770_),
    .X(_03120_));
 sky130_fd_sc_hd__xor2_1 _09714_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__or2_1 _09716_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03121_),
    .X(_03123_));
 sky130_fd_sc_hd__and2_1 _09717_ (.A(_03122_),
    .B(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__inv_2 _09718_ (.A(_03109_),
    .Y(_03125_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__o21a_1 _09720_ (.A1(_03110_),
    .A2(_03115_),
    .B1(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__xnor2_1 _09721_ (.A(_03124_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__or2_1 _09722_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(_03129_));
 sky130_fd_sc_hd__o211a_1 _09723_ (.A1(_02748_),
    .A2(_03128_),
    .B1(_03129_),
    .C1(_03058_),
    .X(_00357_));
 sky130_fd_sc_hd__or3_1 _09724_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .C(_03107_),
    .X(_03130_));
 sky130_fd_sc_hd__and2_1 _09725_ (.A(_02771_),
    .B(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__xnor2_2 _09726_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__xor2_2 _09727_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__a22o_1 _09728_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_03125_),
    .B1(_03121_),
    .B2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(_03134_));
 sky130_fd_sc_hd__or2b_1 _09729_ (.A(_03110_),
    .B_N(_03124_),
    .X(_03135_));
 sky130_fd_sc_hd__nor2_1 _09730_ (.A(_03111_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__nor2_1 _09731_ (.A(_03114_),
    .B(_03135_),
    .Y(_03137_));
 sky130_fd_sc_hd__a221o_2 _09732_ (.A1(_03123_),
    .A2(_03134_),
    .B1(_03136_),
    .B2(_03094_),
    .C1(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__xnor2_1 _09733_ (.A(_03133_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__or2_1 _09734_ (.A(_02804_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_03140_));
 sky130_fd_sc_hd__o211a_1 _09735_ (.A1(_02748_),
    .A2(_03139_),
    .B1(_03140_),
    .C1(_03058_),
    .X(_00358_));
 sky130_fd_sc_hd__o21a_1 _09736_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_03130_),
    .B1(_02772_),
    .X(_03141_));
 sky130_fd_sc_hd__xor2_2 _09737_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__xnor2_1 _09738_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__inv_2 _09739_ (.A(_03132_),
    .Y(_03144_));
 sky130_fd_sc_hd__and2b_1 _09740_ (.A_N(_03133_),
    .B(_03138_),
    .X(_03145_));
 sky130_fd_sc_hd__a21o_1 _09741_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_03144_),
    .B1(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__o21ai_1 _09742_ (.A1(_03143_),
    .A2(_03146_),
    .B1(_02750_),
    .Y(_03147_));
 sky130_fd_sc_hd__a21o_1 _09743_ (.A1(_03143_),
    .A2(_03146_),
    .B1(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__o211a_1 _09744_ (.A1(_02754_),
    .A2(net429),
    .B1(_03017_),
    .C1(_03148_),
    .X(_00359_));
 sky130_fd_sc_hd__nor3_1 _09745_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(_03130_),
    .Y(_03149_));
 sky130_fd_sc_hd__nor2_1 _09746_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__mux2_2 _09747_ (.A0(_03150_),
    .A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .S(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_03151_));
 sky130_fd_sc_hd__a21oi_1 _09748_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A2(_03149_),
    .B1(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__xor2_1 _09749_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__a22o_1 _09750_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_03144_),
    .B1(_03142_),
    .B2(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_03154_));
 sky130_fd_sc_hd__o21ai_1 _09751_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_03142_),
    .B1(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__nor2_1 _09752_ (.A(_03133_),
    .B(_03143_),
    .Y(_03156_));
 sky130_fd_sc_hd__nand2_1 _09753_ (.A(_03138_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__a31o_1 _09754_ (.A1(_03153_),
    .A2(_03155_),
    .A3(_03157_),
    .B1(_02745_),
    .X(_03158_));
 sky130_fd_sc_hd__a21oi_1 _09755_ (.A1(_03155_),
    .A2(_03157_),
    .B1(_03153_),
    .Y(_03159_));
 sky130_fd_sc_hd__a2bb2o_1 _09756_ (.A1_N(_03158_),
    .A2_N(_03159_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B2(_02746_),
    .X(_03160_));
 sky130_fd_sc_hd__and2_1 _09757_ (.A(_03024_),
    .B(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__clkbuf_1 _09758_ (.A(_03161_),
    .X(_00360_));
 sky130_fd_sc_hd__and2b_1 _09759_ (.A_N(_03152_),
    .B(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_03162_));
 sky130_fd_sc_hd__and2_1 _09760_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_03151_),
    .X(_03163_));
 sky130_fd_sc_hd__nor2_1 _09761_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_03151_),
    .Y(_03164_));
 sky130_fd_sc_hd__or2_1 _09762_ (.A(_03163_),
    .B(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__o21a_1 _09763_ (.A1(_03162_),
    .A2(_03159_),
    .B1(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__o31ai_1 _09764_ (.A1(_03162_),
    .A2(_03159_),
    .A3(_03165_),
    .B1(_02751_),
    .Y(_03167_));
 sky130_fd_sc_hd__o221a_1 _09765_ (.A1(_02755_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_03166_),
    .B2(_03167_),
    .C1(_03013_),
    .X(_00361_));
 sky130_fd_sc_hd__and2_1 _09766_ (.A(_02761_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_1 _09767_ (.A(_03153_),
    .B(_03165_),
    .Y(_03169_));
 sky130_fd_sc_hd__and3_1 _09768_ (.A(_03138_),
    .B(_03156_),
    .C(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__o21ba_1 _09769_ (.A1(_03162_),
    .A2(_03163_),
    .B1_N(_03164_),
    .X(_03171_));
 sky130_fd_sc_hd__and2b_1 _09770_ (.A_N(_03155_),
    .B(_03169_),
    .X(_03172_));
 sky130_fd_sc_hd__xor2_1 _09771_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03151_),
    .X(_03173_));
 sky130_fd_sc_hd__o31a_1 _09772_ (.A1(_03170_),
    .A2(_03171_),
    .A3(_03172_),
    .B1(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__or4_1 _09773_ (.A(_03173_),
    .B(_03170_),
    .C(_03171_),
    .D(_03172_),
    .X(_03175_));
 sky130_fd_sc_hd__and3b_1 _09774_ (.A_N(_03174_),
    .B(_03175_),
    .C(_02804_),
    .X(_03176_));
 sky130_fd_sc_hd__o21a_1 _09775_ (.A1(_03168_),
    .A2(_03176_),
    .B1(_02132_),
    .X(_00362_));
 sky130_fd_sc_hd__a21o_1 _09776_ (.A1(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_03151_),
    .B1(_03174_),
    .X(_03177_));
 sky130_fd_sc_hd__xnor2_1 _09777_ (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_03151_),
    .Y(_03178_));
 sky130_fd_sc_hd__xnor2_1 _09778_ (.A(_03177_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__or2_1 _09779_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_02804_),
    .X(_03180_));
 sky130_fd_sc_hd__o211a_1 _09780_ (.A1(_02747_),
    .A2(_03179_),
    .B1(_03180_),
    .C1(_03058_),
    .X(_00363_));
 sky130_fd_sc_hd__and2_1 _09781_ (.A(_02751_),
    .B(_02310_),
    .X(_03181_));
 sky130_fd_sc_hd__clkbuf_1 _09782_ (.A(_03181_),
    .X(_00364_));
 sky130_fd_sc_hd__inv_2 _09783_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_03182_));
 sky130_fd_sc_hd__clkbuf_4 _09784_ (.A(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__buf_4 _09785_ (.A(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_4 _09786_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_4 _09787_ (.A(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__or2_1 _09788_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__o211a_1 _09789_ (.A1(_03184_),
    .A2(net145),
    .B1(_03017_),
    .C1(_03187_),
    .X(_00365_));
 sky130_fd_sc_hd__or2_1 _09790_ (.A(net132),
    .B(_03186_),
    .X(_03188_));
 sky130_fd_sc_hd__o211a_1 _09791_ (.A1(_03184_),
    .A2(net226),
    .B1(_03017_),
    .C1(_03188_),
    .X(_00366_));
 sky130_fd_sc_hd__clkbuf_4 _09792_ (.A(_03186_),
    .X(_03189_));
 sky130_fd_sc_hd__buf_2 _09793_ (.A(_03185_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_4 _09794_ (.A(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__nand2_1 _09795_ (.A(_03191_),
    .B(net305),
    .Y(_03192_));
 sky130_fd_sc_hd__o211a_1 _09796_ (.A1(net141),
    .A2(_03189_),
    .B1(_03017_),
    .C1(_03192_),
    .X(_00367_));
 sky130_fd_sc_hd__or2_1 _09797_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_03193_));
 sky130_fd_sc_hd__nand2_1 _09798_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .Y(_03194_));
 sky130_fd_sc_hd__and3_1 _09799_ (.A(_02851_),
    .B(_03193_),
    .C(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__a21oi_1 _09800_ (.A1(_03193_),
    .A2(_03194_),
    .B1(_02851_),
    .Y(_03196_));
 sky130_fd_sc_hd__o21ai_1 _09801_ (.A1(_03195_),
    .A2(_03196_),
    .B1(_03191_),
    .Y(_03197_));
 sky130_fd_sc_hd__o211a_1 _09802_ (.A1(net136),
    .A2(_03189_),
    .B1(_03017_),
    .C1(_03197_),
    .X(_00368_));
 sky130_fd_sc_hd__or2_1 _09803_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(_03193_),
    .X(_03198_));
 sky130_fd_sc_hd__nand2_1 _09804_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(_03193_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_1 _09805_ (.A1(_03198_),
    .A2(_03199_),
    .B1(_03196_),
    .Y(_03200_));
 sky130_fd_sc_hd__clkbuf_4 _09806_ (.A(_03182_),
    .X(_03201_));
 sky130_fd_sc_hd__a31o_1 _09807_ (.A1(_03196_),
    .A2(_03198_),
    .A3(_03199_),
    .B1(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__o221a_1 _09808_ (.A1(net130),
    .A2(_03189_),
    .B1(_03200_),
    .B2(_03202_),
    .C1(_03013_),
    .X(_00369_));
 sky130_fd_sc_hd__inv_2 _09809_ (.A(_03198_),
    .Y(_03203_));
 sky130_fd_sc_hd__and3_1 _09810_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .C(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_03204_));
 sky130_fd_sc_hd__inv_2 _09811_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_03205_));
 sky130_fd_sc_hd__buf_2 _09812_ (.A(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_4 _09813_ (.A(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__mux2_1 _09814_ (.A0(_03203_),
    .A1(_03204_),
    .S(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__xnor2_1 _09815_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_1 _09816_ (.A(_03191_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__o211a_1 _09817_ (.A1(net266),
    .A2(_03189_),
    .B1(_03017_),
    .C1(_03210_),
    .X(_00370_));
 sky130_fd_sc_hd__nand2_1 _09818_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_03204_),
    .Y(_03211_));
 sky130_fd_sc_hd__or2_1 _09819_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_03198_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_1 _09820_ (.A0(_03211_),
    .A1(_03212_),
    .S(_02850_),
    .X(_03213_));
 sky130_fd_sc_hd__xnor2_1 _09821_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__or2_1 _09822_ (.A(net254),
    .B(_03190_),
    .X(_03215_));
 sky130_fd_sc_hd__o211a_1 _09823_ (.A1(_03184_),
    .A2(net496),
    .B1(_03215_),
    .C1(_03058_),
    .X(_00371_));
 sky130_fd_sc_hd__or2_1 _09824_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_03212_),
    .X(_03216_));
 sky130_fd_sc_hd__a31o_1 _09825_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A3(_03204_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_03217_));
 sky130_fd_sc_hd__a21bo_1 _09826_ (.A1(_02851_),
    .A2(_03216_),
    .B1_N(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__xnor2_1 _09827_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__or2_1 _09828_ (.A(net126),
    .B(_03190_),
    .X(_03220_));
 sky130_fd_sc_hd__o211a_1 _09829_ (.A1(_03184_),
    .A2(_03219_),
    .B1(_03220_),
    .C1(_03058_),
    .X(_00372_));
 sky130_fd_sc_hd__and4_1 _09830_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .D(_03204_),
    .X(_03221_));
 sky130_fd_sc_hd__o21ai_1 _09831_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(_03216_),
    .B1(_02851_),
    .Y(_03222_));
 sky130_fd_sc_hd__o21ai_1 _09832_ (.A1(_02851_),
    .A2(_03221_),
    .B1(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__xnor2_1 _09833_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__or2_1 _09834_ (.A(net124),
    .B(_03190_),
    .X(_03225_));
 sky130_fd_sc_hd__o211a_1 _09835_ (.A1(_03184_),
    .A2(_03224_),
    .B1(_03225_),
    .C1(_03058_),
    .X(_00373_));
 sky130_fd_sc_hd__or3_1 _09836_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .C(_03216_),
    .X(_03226_));
 sky130_fd_sc_hd__or2_1 _09837_ (.A(_03207_),
    .B(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__and2_1 _09838_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_03221_),
    .X(_03228_));
 sky130_fd_sc_hd__nand2_1 _09839_ (.A(_03207_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21oi_1 _09840_ (.A1(_03227_),
    .A2(_03229_),
    .B1(net395),
    .Y(_03230_));
 sky130_fd_sc_hd__a31o_1 _09841_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(_03227_),
    .A3(_03229_),
    .B1(_03201_),
    .X(_03231_));
 sky130_fd_sc_hd__o221a_1 _09842_ (.A1(net298),
    .A2(_03189_),
    .B1(_03230_),
    .B2(_03231_),
    .C1(_03013_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _09843_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_03228_),
    .Y(_03232_));
 sky130_fd_sc_hd__or2_1 _09844_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_03226_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(_03232_),
    .A1(_03233_),
    .S(_02850_),
    .X(_03234_));
 sky130_fd_sc_hd__nor2_1 _09846_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__a21o_1 _09847_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_03234_),
    .B1(_03183_),
    .X(_03236_));
 sky130_fd_sc_hd__o221a_1 _09848_ (.A1(net252),
    .A2(_03189_),
    .B1(_03235_),
    .B2(_03236_),
    .C1(_03013_),
    .X(_00375_));
 sky130_fd_sc_hd__clkbuf_4 _09849_ (.A(_03190_),
    .X(_03237_));
 sky130_fd_sc_hd__or2_1 _09850_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_03233_),
    .X(_03238_));
 sky130_fd_sc_hd__a31o_1 _09851_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A3(_03228_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_03239_));
 sky130_fd_sc_hd__a21bo_1 _09852_ (.A1(_02851_),
    .A2(_03238_),
    .B1_N(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__nor2_1 _09853_ (.A(net580),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__a21o_1 _09854_ (.A1(net603),
    .A2(_03240_),
    .B1(_03183_),
    .X(_03242_));
 sky130_fd_sc_hd__o221a_1 _09855_ (.A1(_03237_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_03241_),
    .B2(_03242_),
    .C1(_03013_),
    .X(_00376_));
 sky130_fd_sc_hd__and4_1 _09856_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .D(_03228_),
    .X(_03243_));
 sky130_fd_sc_hd__or2_1 _09857_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_03238_),
    .X(_03244_));
 sky130_fd_sc_hd__inv_2 _09858_ (.A(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__mux2_1 _09859_ (.A0(_03243_),
    .A1(_03245_),
    .S(_02850_),
    .X(_03246_));
 sky130_fd_sc_hd__nor2_1 _09860_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__a21o_1 _09861_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_03246_),
    .B1(_03183_),
    .X(_03248_));
 sky130_fd_sc_hd__o221a_1 _09862_ (.A1(_03237_),
    .A2(net487),
    .B1(_03247_),
    .B2(_03248_),
    .C1(_03013_),
    .X(_00377_));
 sky130_fd_sc_hd__or3_1 _09863_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_03243_),
    .X(_03249_));
 sky130_fd_sc_hd__o21ai_1 _09864_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_03243_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .Y(_03250_));
 sky130_fd_sc_hd__a21oi_1 _09865_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_02851_),
    .Y(_03251_));
 sky130_fd_sc_hd__a21o_1 _09866_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_03244_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(_03252_));
 sky130_fd_sc_hd__nand3_2 _09867_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_03244_),
    .Y(_03253_));
 sky130_fd_sc_hd__a31o_1 _09868_ (.A1(_02851_),
    .A2(_03252_),
    .A3(_03253_),
    .B1(_03201_),
    .X(_03254_));
 sky130_fd_sc_hd__o221a_1 _09869_ (.A1(_03237_),
    .A2(net532),
    .B1(_03251_),
    .B2(_03254_),
    .C1(_03013_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _09870_ (.A0(_03249_),
    .A1(_03253_),
    .S(_02850_),
    .X(_03255_));
 sky130_fd_sc_hd__nor2_1 _09871_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__a21o_1 _09872_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_03255_),
    .B1(_03183_),
    .X(_03257_));
 sky130_fd_sc_hd__clkbuf_4 _09873_ (.A(_02308_),
    .X(_03258_));
 sky130_fd_sc_hd__o221a_1 _09874_ (.A1(_03237_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_03256_),
    .B2(_03257_),
    .C1(_03258_),
    .X(_00379_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(_02850_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .Y(_03259_));
 sky130_fd_sc_hd__or2_1 _09876_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_03249_),
    .X(_03260_));
 sky130_fd_sc_hd__o22a_1 _09877_ (.A1(_03253_),
    .A2(_03259_),
    .B1(_03260_),
    .B2(_02850_),
    .X(_03261_));
 sky130_fd_sc_hd__and2_1 _09878_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__o21ai_1 _09879_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_03261_),
    .B1(_03186_),
    .Y(_03263_));
 sky130_fd_sc_hd__o221a_1 _09880_ (.A1(_03237_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_03262_),
    .B2(_03263_),
    .C1(_03258_),
    .X(_00380_));
 sky130_fd_sc_hd__inv_2 _09881_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .Y(_03264_));
 sky130_fd_sc_hd__nor2_1 _09882_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_03260_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _09883_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .Y(_03266_));
 sky130_fd_sc_hd__o21ai_1 _09884_ (.A1(_03253_),
    .A2(_03266_),
    .B1(_02850_),
    .Y(_03267_));
 sky130_fd_sc_hd__o21a_1 _09885_ (.A1(_02851_),
    .A2(_03265_),
    .B1(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__nor2_1 _09886_ (.A(_03264_),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__a21o_1 _09887_ (.A1(_03264_),
    .A2(_03268_),
    .B1(_03183_),
    .X(_03270_));
 sky130_fd_sc_hd__o221a_1 _09888_ (.A1(_03237_),
    .A2(net541),
    .B1(_03269_),
    .B2(_03270_),
    .C1(_03258_),
    .X(_00381_));
 sky130_fd_sc_hd__inv_2 _09889_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .Y(_03271_));
 sky130_fd_sc_hd__a21o_1 _09890_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_02850_),
    .X(_03272_));
 sky130_fd_sc_hd__o211a_1 _09891_ (.A1(_03207_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_03267_),
    .C1(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__xnor2_1 _09892_ (.A(_03271_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__or2_1 _09893_ (.A(_03186_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(_03275_));
 sky130_fd_sc_hd__o211a_1 _09894_ (.A1(_03184_),
    .A2(_03274_),
    .B1(_03275_),
    .C1(_03058_),
    .X(_00382_));
 sky130_fd_sc_hd__o41a_1 _09895_ (.A1(_03271_),
    .A2(_03264_),
    .A3(_03253_),
    .A4(_03266_),
    .B1(_02850_),
    .X(_03276_));
 sky130_fd_sc_hd__o41a_1 _09896_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A4(_03260_),
    .B1(_03207_),
    .X(_03277_));
 sky130_fd_sc_hd__o21a_1 _09897_ (.A1(_03276_),
    .A2(_03277_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_03278_));
 sky130_fd_sc_hd__o31ai_1 _09898_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_03276_),
    .A3(_03277_),
    .B1(_03186_),
    .Y(_03279_));
 sky130_fd_sc_hd__o221a_1 _09899_ (.A1(_03237_),
    .A2(net526),
    .B1(_03278_),
    .B2(_03279_),
    .C1(_03258_),
    .X(_00383_));
 sky130_fd_sc_hd__clkbuf_4 _09900_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_03280_));
 sky130_fd_sc_hd__and2b_1 _09901_ (.A_N(_03276_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_03281_));
 sky130_fd_sc_hd__o21ai_1 _09902_ (.A1(_03277_),
    .A2(_03281_),
    .B1(_03191_),
    .Y(_03282_));
 sky130_fd_sc_hd__o211a_1 _09903_ (.A1(_03189_),
    .A2(_03280_),
    .B1(_03017_),
    .C1(_03282_),
    .X(_00384_));
 sky130_fd_sc_hd__inv_2 _09904_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_03283_));
 sky130_fd_sc_hd__nor2_1 _09905_ (.A(_03283_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_03284_));
 sky130_fd_sc_hd__a21o_1 _09906_ (.A1(_03283_),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_03183_),
    .X(_03285_));
 sky130_fd_sc_hd__o221a_1 _09907_ (.A1(_03237_),
    .A2(net431),
    .B1(_03284_),
    .B2(_03285_),
    .C1(_03258_),
    .X(_00385_));
 sky130_fd_sc_hd__and2b_1 _09908_ (.A_N(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_03286_));
 sky130_fd_sc_hd__xnor2_1 _09909_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__xnor2_1 _09910_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__xor2_1 _09911_ (.A(_03284_),
    .B(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__buf_2 _09912_ (.A(_03185_),
    .X(_03290_));
 sky130_fd_sc_hd__or2_1 _09913_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_03291_));
 sky130_fd_sc_hd__clkbuf_4 _09914_ (.A(_01474_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_1 _09915_ (.A1(_03184_),
    .A2(_03289_),
    .B1(_03291_),
    .C1(_03292_),
    .X(_00386_));
 sky130_fd_sc_hd__and2_1 _09916_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_03287_),
    .X(_03293_));
 sky130_fd_sc_hd__nor2_1 _09917_ (.A(_03284_),
    .B(_03288_),
    .Y(_03294_));
 sky130_fd_sc_hd__o21ba_1 _09918_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B1_N(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_03295_));
 sky130_fd_sc_hd__xnor2_1 _09919_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__or2_1 _09920_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_03296_),
    .Y(_03298_));
 sky130_fd_sc_hd__and2_1 _09922_ (.A(_03297_),
    .B(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o21ai_1 _09923_ (.A1(_03293_),
    .A2(_03294_),
    .B1(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__o31a_1 _09924_ (.A1(_03293_),
    .A2(_03294_),
    .A3(_03299_),
    .B1(_03185_),
    .X(_03301_));
 sky130_fd_sc_hd__a22oi_1 _09925_ (.A1(_03201_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_03300_),
    .B2(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__and2b_1 _09926_ (.A_N(_03302_),
    .B(_03118_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _09927_ (.A(_03303_),
    .X(_00387_));
 sky130_fd_sc_hd__o31a_1 _09928_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A3(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B1(_03205_),
    .X(_03304_));
 sky130_fd_sc_hd__xnor2_1 _09929_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__and2_1 _09930_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__nor2_1 _09931_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_03305_),
    .Y(_03307_));
 sky130_fd_sc_hd__or2_1 _09932_ (.A(_03306_),
    .B(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__and3_1 _09933_ (.A(_03298_),
    .B(_03300_),
    .C(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__a21oi_1 _09934_ (.A1(_03298_),
    .A2(_03300_),
    .B1(_03308_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_1 _09935_ (.A(_03182_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .Y(_03311_));
 sky130_fd_sc_hd__o31a_1 _09936_ (.A1(_03182_),
    .A2(_03309_),
    .A3(_03310_),
    .B1(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__and2b_1 _09937_ (.A_N(_03312_),
    .B(_03118_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _09938_ (.A(_03313_),
    .X(_00388_));
 sky130_fd_sc_hd__or2_1 _09939_ (.A(_03306_),
    .B(_03310_),
    .X(_03314_));
 sky130_fd_sc_hd__or4_4 _09940_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .C(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .D(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_03315_));
 sky130_fd_sc_hd__nand2_1 _09941_ (.A(_03205_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__xor2_1 _09942_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__and2_1 _09943_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__nor2_1 _09944_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_03317_),
    .Y(_03319_));
 sky130_fd_sc_hd__nor2_1 _09945_ (.A(_03318_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__xor2_1 _09946_ (.A(_03314_),
    .B(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__or2_1 _09947_ (.A(_03290_),
    .B(net614),
    .X(_03322_));
 sky130_fd_sc_hd__o211a_1 _09948_ (.A1(_03184_),
    .A2(_03321_),
    .B1(_03322_),
    .C1(_03292_),
    .X(_00389_));
 sky130_fd_sc_hd__o21a_1 _09949_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_03315_),
    .B1(_03205_),
    .X(_03323_));
 sky130_fd_sc_hd__xor2_1 _09950_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__and2b_1 _09951_ (.A_N(_03324_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_03325_));
 sky130_fd_sc_hd__or2b_1 _09952_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B_N(_03324_),
    .X(_03326_));
 sky130_fd_sc_hd__and2b_1 _09953_ (.A_N(_03325_),
    .B(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__a21o_1 _09954_ (.A1(_03314_),
    .A2(_03320_),
    .B1(_03318_),
    .X(_03328_));
 sky130_fd_sc_hd__xnor2_1 _09955_ (.A(_03327_),
    .B(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _09956_ (.A(_03191_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__o211a_1 _09957_ (.A1(_03189_),
    .A2(net441),
    .B1(_03017_),
    .C1(_03330_),
    .X(_00390_));
 sky130_fd_sc_hd__o31a_1 _09958_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A3(_03315_),
    .B1(_03205_),
    .X(_03331_));
 sky130_fd_sc_hd__xnor2_1 _09959_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__and2_1 _09960_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__nor2_1 _09961_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03332_),
    .Y(_03334_));
 sky130_fd_sc_hd__nor2_1 _09962_ (.A(_03333_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__and2_1 _09963_ (.A(_03320_),
    .B(_03327_),
    .X(_03336_));
 sky130_fd_sc_hd__o21a_1 _09964_ (.A1(_03318_),
    .A2(_03325_),
    .B1(_03326_),
    .X(_03337_));
 sky130_fd_sc_hd__a21oi_1 _09965_ (.A1(_03314_),
    .A2(_03336_),
    .B1(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__xnor2_1 _09966_ (.A(_03335_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A1(_03339_),
    .S(_03185_),
    .X(_03340_));
 sky130_fd_sc_hd__and2_1 _09968_ (.A(_03024_),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_1 _09969_ (.A(_03341_),
    .X(_00391_));
 sky130_fd_sc_hd__a21o_1 _09970_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_03205_),
    .B1(_03331_),
    .X(_03342_));
 sky130_fd_sc_hd__xor2_1 _09971_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__or2b_1 _09972_ (.A(_03343_),
    .B_N(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_03344_));
 sky130_fd_sc_hd__or2b_1 _09973_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B_N(_03343_),
    .X(_03345_));
 sky130_fd_sc_hd__and2_1 _09974_ (.A(_03344_),
    .B(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03332_),
    .Y(_03347_));
 sky130_fd_sc_hd__o21ai_1 _09976_ (.A1(_03334_),
    .A2(_03338_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__xor2_1 _09977_ (.A(_03346_),
    .B(_03348_),
    .X(_03349_));
 sky130_fd_sc_hd__or2_1 _09978_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_03350_));
 sky130_fd_sc_hd__o211a_1 _09979_ (.A1(_03184_),
    .A2(_03349_),
    .B1(_03350_),
    .C1(_03292_),
    .X(_00392_));
 sky130_fd_sc_hd__nand2_1 _09980_ (.A(_03347_),
    .B(_03344_),
    .Y(_03351_));
 sky130_fd_sc_hd__a32o_1 _09981_ (.A1(_03335_),
    .A2(_03337_),
    .A3(_03346_),
    .B1(_03351_),
    .B2(_03345_),
    .X(_03352_));
 sky130_fd_sc_hd__o2111a_1 _09982_ (.A1(_03306_),
    .A2(_03310_),
    .B1(_03335_),
    .C1(_03336_),
    .D1(_03346_),
    .X(_03353_));
 sky130_fd_sc_hd__nor2_1 _09983_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__or2_1 _09984_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .X(_03355_));
 sky130_fd_sc_hd__or4_4 _09985_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .C(_03315_),
    .D(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__and2_1 _09986_ (.A(_03206_),
    .B(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__xnor2_1 _09987_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__nand2_1 _09988_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__or2_1 _09989_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03358_),
    .X(_03360_));
 sky130_fd_sc_hd__nand2_1 _09990_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xor2_1 _09991_ (.A(_03354_),
    .B(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__or2_1 _09992_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_03363_));
 sky130_fd_sc_hd__o211a_1 _09993_ (.A1(_03184_),
    .A2(_03362_),
    .B1(_03363_),
    .C1(_03292_),
    .X(_00393_));
 sky130_fd_sc_hd__o21bai_2 _09994_ (.A1(_03352_),
    .A2(_03353_),
    .B1_N(_03361_),
    .Y(_03364_));
 sky130_fd_sc_hd__o21a_1 _09995_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_03356_),
    .B1(_03206_),
    .X(_03365_));
 sky130_fd_sc_hd__xor2_2 _09996_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__xnor2_2 _09997_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__a21oi_1 _09998_ (.A1(_03359_),
    .A2(_03364_),
    .B1(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__a31o_1 _09999_ (.A1(_03359_),
    .A2(_03364_),
    .A3(_03367_),
    .B1(_03201_),
    .X(_03369_));
 sky130_fd_sc_hd__o221a_1 _10000_ (.A1(_03237_),
    .A2(net550),
    .B1(_03368_),
    .B2(_03369_),
    .C1(_03258_),
    .X(_00394_));
 sky130_fd_sc_hd__or3_2 _10001_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .C(_03356_),
    .X(_03370_));
 sky130_fd_sc_hd__and2_1 _10002_ (.A(_03206_),
    .B(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__xnor2_1 _10003_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__xor2_1 _10004_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__inv_2 _10005_ (.A(_03367_),
    .Y(_03374_));
 sky130_fd_sc_hd__inv_2 _10006_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .Y(_03375_));
 sky130_fd_sc_hd__o21a_1 _10007_ (.A1(_03375_),
    .A2(_03366_),
    .B1(_03359_),
    .X(_03376_));
 sky130_fd_sc_hd__a21o_1 _10008_ (.A1(_03375_),
    .A2(_03366_),
    .B1(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__o21ai_1 _10009_ (.A1(_03364_),
    .A2(_03374_),
    .B1(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__nand2_1 _10010_ (.A(_03373_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__o21a_1 _10011_ (.A1(_03373_),
    .A2(_03378_),
    .B1(_03185_),
    .X(_03380_));
 sky130_fd_sc_hd__a22o_1 _10012_ (.A1(_03201_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_03379_),
    .B2(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__and2_1 _10013_ (.A(_03024_),
    .B(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_1 _10014_ (.A(_03382_),
    .X(_00395_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03372_),
    .Y(_03383_));
 sky130_fd_sc_hd__o21a_1 _10016_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_03370_),
    .B1(_03206_),
    .X(_03384_));
 sky130_fd_sc_hd__xor2_1 _10017_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__xnor2_1 _10018_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__a21oi_1 _10019_ (.A1(_03383_),
    .A2(_03379_),
    .B1(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a31o_1 _10020_ (.A1(_03383_),
    .A2(_03379_),
    .A3(_03386_),
    .B1(_03201_),
    .X(_03388_));
 sky130_fd_sc_hd__o221a_1 _10021_ (.A1(_03191_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_03387_),
    .B2(_03388_),
    .C1(_03258_),
    .X(_00396_));
 sky130_fd_sc_hd__clkbuf_4 _10022_ (.A(_03183_),
    .X(_03389_));
 sky130_fd_sc_hd__or2_1 _10023_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_03390_));
 sky130_fd_sc_hd__or2_1 _10024_ (.A(_03370_),
    .B(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__and2_1 _10025_ (.A(_03207_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__xnor2_1 _10026_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__and2_1 _10027_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__nor2_1 _10028_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_03393_),
    .Y(_03395_));
 sky130_fd_sc_hd__or2_1 _10029_ (.A(_03394_),
    .B(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__nand2_1 _10030_ (.A(_03373_),
    .B(_03386_),
    .Y(_03397_));
 sky130_fd_sc_hd__inv_2 _10031_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .Y(_03398_));
 sky130_fd_sc_hd__o21a_1 _10032_ (.A1(_03398_),
    .A2(_03385_),
    .B1(_03383_),
    .X(_03399_));
 sky130_fd_sc_hd__and2_1 _10033_ (.A(_03398_),
    .B(_03385_),
    .X(_03400_));
 sky130_fd_sc_hd__o22a_1 _10034_ (.A1(_03377_),
    .A2(_03397_),
    .B1(_03399_),
    .B2(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__o31a_1 _10035_ (.A1(_03364_),
    .A2(_03374_),
    .A3(_03397_),
    .B1(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__or2_1 _10036_ (.A(_03396_),
    .B(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(_03396_),
    .B(_03402_),
    .Y(_03404_));
 sky130_fd_sc_hd__and2_1 _10038_ (.A(_03403_),
    .B(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__or2_1 _10039_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_03406_));
 sky130_fd_sc_hd__o211a_1 _10040_ (.A1(_03389_),
    .A2(_03405_),
    .B1(_03406_),
    .C1(_03292_),
    .X(_00397_));
 sky130_fd_sc_hd__inv_2 _10041_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_03407_));
 sky130_fd_sc_hd__o21ai_1 _10042_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_03391_),
    .B1(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__mux2_1 _10043_ (.A0(_03407_),
    .A1(_03408_),
    .S(_03207_),
    .X(_03409_));
 sky130_fd_sc_hd__buf_2 _10044_ (.A(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__or3_1 _10045_ (.A(_03407_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .C(_03391_),
    .X(_03411_));
 sky130_fd_sc_hd__a21oi_1 _10046_ (.A1(_03410_),
    .A2(_03411_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .Y(_03412_));
 sky130_fd_sc_hd__and3_1 _10047_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_03410_),
    .C(_03411_),
    .X(_03413_));
 sky130_fd_sc_hd__nor2_1 _10048_ (.A(_03412_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__and2b_1 _10049_ (.A_N(_03394_),
    .B(_03403_),
    .X(_03415_));
 sky130_fd_sc_hd__and2_1 _10050_ (.A(_03414_),
    .B(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__o21ai_1 _10051_ (.A1(_03414_),
    .A2(_03415_),
    .B1(_03186_),
    .Y(_03417_));
 sky130_fd_sc_hd__o221a_1 _10052_ (.A1(_03191_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_03416_),
    .B2(_03417_),
    .C1(_03258_),
    .X(_00398_));
 sky130_fd_sc_hd__nand2_1 _10053_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03410_),
    .Y(_03418_));
 sky130_fd_sc_hd__or2_1 _10054_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03410_),
    .X(_03419_));
 sky130_fd_sc_hd__and2_1 _10055_ (.A(_03418_),
    .B(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__nor2_1 _10056_ (.A(_03394_),
    .B(_03413_),
    .Y(_03421_));
 sky130_fd_sc_hd__a21o_1 _10057_ (.A1(_03403_),
    .A2(_03421_),
    .B1(_03412_),
    .X(_03422_));
 sky130_fd_sc_hd__xnor2_1 _10058_ (.A(_03420_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__mux2_1 _10059_ (.A0(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A1(_03423_),
    .S(_03185_),
    .X(_03424_));
 sky130_fd_sc_hd__and2_1 _10060_ (.A(_03024_),
    .B(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__clkbuf_1 _10061_ (.A(_03425_),
    .X(_00399_));
 sky130_fd_sc_hd__xor2_1 _10062_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_03410_),
    .X(_03426_));
 sky130_fd_sc_hd__inv_2 _10063_ (.A(_03420_),
    .Y(_03427_));
 sky130_fd_sc_hd__o21ai_1 _10064_ (.A1(_03427_),
    .A2(_03422_),
    .B1(_03418_),
    .Y(_03428_));
 sky130_fd_sc_hd__xor2_1 _10065_ (.A(_03426_),
    .B(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__or2_1 _10066_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(_03430_));
 sky130_fd_sc_hd__o211a_1 _10067_ (.A1(_03389_),
    .A2(_03429_),
    .B1(_03430_),
    .C1(_03292_),
    .X(_00400_));
 sky130_fd_sc_hd__nor2_1 _10068_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03410_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _10069_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03410_),
    .Y(_03432_));
 sky130_fd_sc_hd__and2b_1 _10070_ (.A_N(_03431_),
    .B(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__and2_1 _10071_ (.A(_03420_),
    .B(_03426_),
    .X(_03434_));
 sky130_fd_sc_hd__nand2_1 _10072_ (.A(_03414_),
    .B(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__or3b_1 _10073_ (.A(_03412_),
    .B(_03421_),
    .C_N(_03434_),
    .X(_03436_));
 sky130_fd_sc_hd__o21ai_1 _10074_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_03410_),
    .Y(_03437_));
 sky130_fd_sc_hd__o211a_1 _10075_ (.A1(_03403_),
    .A2(_03435_),
    .B1(_03436_),
    .C1(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__xnor2_1 _10076_ (.A(_03433_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__mux2_1 _10077_ (.A0(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A1(_03439_),
    .S(_03185_),
    .X(_03440_));
 sky130_fd_sc_hd__and2_1 _10078_ (.A(_03024_),
    .B(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_1 _10079_ (.A(_03441_),
    .X(_00401_));
 sky130_fd_sc_hd__o21ai_1 _10080_ (.A1(_03431_),
    .A2(_03438_),
    .B1(_03432_),
    .Y(_03442_));
 sky130_fd_sc_hd__xnor2_1 _10081_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_03410_),
    .Y(_03443_));
 sky130_fd_sc_hd__xnor2_1 _10082_ (.A(_03442_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__or2_1 _10083_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_03445_));
 sky130_fd_sc_hd__o211a_1 _10084_ (.A1(_03389_),
    .A2(_03444_),
    .B1(_03445_),
    .C1(_03292_),
    .X(_00402_));
 sky130_fd_sc_hd__and2_1 _10085_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(_03446_));
 sky130_fd_sc_hd__nor2_1 _10086_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .Y(_03447_));
 sky130_fd_sc_hd__o21ai_1 _10087_ (.A1(_03446_),
    .A2(_03447_),
    .B1(_03191_),
    .Y(_03448_));
 sky130_fd_sc_hd__o211a_1 _10088_ (.A1(_03189_),
    .A2(net297),
    .B1(_03017_),
    .C1(_03448_),
    .X(_00403_));
 sky130_fd_sc_hd__and2b_1 _10089_ (.A_N(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(_03449_));
 sky130_fd_sc_hd__xnor2_1 _10090_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__xnor2_1 _10091_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__xor2_1 _10092_ (.A(_03446_),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__or2_1 _10093_ (.A(_03290_),
    .B(net620),
    .X(_03453_));
 sky130_fd_sc_hd__o211a_1 _10094_ (.A1(_03389_),
    .A2(_03452_),
    .B1(_03453_),
    .C1(_03292_),
    .X(_00404_));
 sky130_fd_sc_hd__o21a_1 _10095_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B1(_03205_),
    .X(_03454_));
 sky130_fd_sc_hd__xnor2_1 _10096_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__and2_1 _10097_ (.A(_03031_),
    .B(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__nor2_1 _10098_ (.A(_03031_),
    .B(_03455_),
    .Y(_03457_));
 sky130_fd_sc_hd__nor2_1 _10099_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__and2b_1 _10100_ (.A_N(_03450_),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_03459_));
 sky130_fd_sc_hd__a21o_1 _10101_ (.A1(_03446_),
    .A2(_03451_),
    .B1(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__nand2_1 _10102_ (.A(_03458_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__o21a_1 _10103_ (.A1(_03458_),
    .A2(_03460_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03462_));
 sky130_fd_sc_hd__a22o_1 _10104_ (.A1(_03182_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_03461_),
    .B2(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__and2_1 _10105_ (.A(_03024_),
    .B(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_1 _10106_ (.A(_03464_),
    .X(_00405_));
 sky130_fd_sc_hd__o31a_1 _10107_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A3(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B1(_03206_),
    .X(_03465_));
 sky130_fd_sc_hd__xnor2_1 _10108_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__nor2_1 _10109_ (.A(_03035_),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand2_1 _10110_ (.A(_03035_),
    .B(_03466_),
    .Y(_03468_));
 sky130_fd_sc_hd__and2b_1 _10111_ (.A_N(_03467_),
    .B(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(_03031_),
    .B(_03455_),
    .Y(_03470_));
 sky130_fd_sc_hd__a21o_1 _10113_ (.A1(_03470_),
    .A2(_03460_),
    .B1(_03457_),
    .X(_03471_));
 sky130_fd_sc_hd__a21o_1 _10114_ (.A1(_03469_),
    .A2(_03471_),
    .B1(_03182_),
    .X(_03472_));
 sky130_fd_sc_hd__nor2_1 _10115_ (.A(_03469_),
    .B(_03471_),
    .Y(_03473_));
 sky130_fd_sc_hd__a2bb2o_1 _10116_ (.A1_N(_03472_),
    .A2_N(_03473_),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B2(_03182_),
    .X(_03474_));
 sky130_fd_sc_hd__and2_1 _10117_ (.A(_03024_),
    .B(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _10118_ (.A(_03475_),
    .X(_00406_));
 sky130_fd_sc_hd__a21oi_2 _10119_ (.A1(_03468_),
    .A2(_03471_),
    .B1(_03467_),
    .Y(_03476_));
 sky130_fd_sc_hd__or4_2 _10120_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .C(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .D(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(_03477_));
 sky130_fd_sc_hd__nand2_1 _10121_ (.A(_03205_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__xor2_1 _10122_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__or2_1 _10123_ (.A(_03283_),
    .B(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__nand2_1 _10124_ (.A(_03283_),
    .B(_03479_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2_1 _10125_ (.A(_03480_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__xor2_1 _10126_ (.A(_03476_),
    .B(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__or2_1 _10127_ (.A(_03290_),
    .B(net503),
    .X(_03484_));
 sky130_fd_sc_hd__o211a_1 _10128_ (.A1(_03389_),
    .A2(_03483_),
    .B1(_03484_),
    .C1(_03292_),
    .X(_00407_));
 sky130_fd_sc_hd__o21a_1 _10129_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_03477_),
    .B1(_03205_),
    .X(_03485_));
 sky130_fd_sc_hd__xnor2_1 _10130_ (.A(_03375_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _10131_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__inv_2 _10132_ (.A(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__nor2_1 _10133_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03486_),
    .Y(_03489_));
 sky130_fd_sc_hd__nor2_1 _10134_ (.A(_03488_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__o21a_1 _10135_ (.A1(_03476_),
    .A2(_03482_),
    .B1(_03480_),
    .X(_03491_));
 sky130_fd_sc_hd__xnor2_1 _10136_ (.A(_03490_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__or2_1 _10137_ (.A(_03290_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_03493_));
 sky130_fd_sc_hd__o211a_1 _10138_ (.A1(_03389_),
    .A2(_03492_),
    .B1(_03493_),
    .C1(_03292_),
    .X(_00408_));
 sky130_fd_sc_hd__inv_2 _10139_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_03494_));
 sky130_fd_sc_hd__o31a_1 _10140_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A3(_03477_),
    .B1(_03205_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_1 _10141_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__nor2_1 _10142_ (.A(_03494_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__nand2_1 _10143_ (.A(_03494_),
    .B(_03496_),
    .Y(_03498_));
 sky130_fd_sc_hd__or2b_1 _10144_ (.A(_03497_),
    .B_N(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__or3_1 _10145_ (.A(_03482_),
    .B(_03488_),
    .C(_03489_),
    .X(_03500_));
 sky130_fd_sc_hd__a21oi_1 _10146_ (.A1(_03480_),
    .A2(_03487_),
    .B1(_03489_),
    .Y(_03501_));
 sky130_fd_sc_hd__inv_2 _10147_ (.A(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__o21ai_1 _10148_ (.A1(_03476_),
    .A2(_03500_),
    .B1(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__xnor2_1 _10149_ (.A(_03499_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_03504_),
    .S(_03185_),
    .X(_03505_));
 sky130_fd_sc_hd__and2_1 _10151_ (.A(_03024_),
    .B(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _10152_ (.A(_03506_),
    .X(_00409_));
 sky130_fd_sc_hd__a21o_1 _10153_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_03206_),
    .B1(_03495_),
    .X(_03507_));
 sky130_fd_sc_hd__xnor2_1 _10154_ (.A(_03398_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__and2_1 _10155_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__nor2_1 _10156_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03508_),
    .Y(_03510_));
 sky130_fd_sc_hd__or2_1 _10157_ (.A(_03509_),
    .B(_03510_),
    .X(_03511_));
 sky130_fd_sc_hd__a21oi_1 _10158_ (.A1(_03498_),
    .A2(_03503_),
    .B1(_03497_),
    .Y(_03512_));
 sky130_fd_sc_hd__xor2_1 _10159_ (.A(_03511_),
    .B(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__or2_1 _10160_ (.A(_03190_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_03514_));
 sky130_fd_sc_hd__buf_4 _10161_ (.A(_01474_),
    .X(_03515_));
 sky130_fd_sc_hd__o211a_1 _10162_ (.A1(_03389_),
    .A2(_03513_),
    .B1(_03514_),
    .C1(_03515_),
    .X(_00410_));
 sky130_fd_sc_hd__nor2_1 _10163_ (.A(_03497_),
    .B(_03509_),
    .Y(_03516_));
 sky130_fd_sc_hd__o32a_1 _10164_ (.A1(_03499_),
    .A2(_03502_),
    .A3(_03511_),
    .B1(_03516_),
    .B2(_03510_),
    .X(_03517_));
 sky130_fd_sc_hd__or4_1 _10165_ (.A(_03476_),
    .B(_03499_),
    .C(_03500_),
    .D(_03511_),
    .X(_03518_));
 sky130_fd_sc_hd__and2_1 _10166_ (.A(_03517_),
    .B(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__or2_1 _10167_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_03520_));
 sky130_fd_sc_hd__or4_4 _10168_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .C(_03477_),
    .D(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__nand2_1 _10169_ (.A(_03206_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__xnor2_1 _10170_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__or2_1 _10172_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_03523_),
    .X(_03525_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(_03524_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__xor2_1 _10174_ (.A(_03519_),
    .B(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__or2_1 _10175_ (.A(_03190_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_03528_));
 sky130_fd_sc_hd__o211a_1 _10176_ (.A1(_03389_),
    .A2(_03527_),
    .B1(_03528_),
    .C1(_03515_),
    .X(_00411_));
 sky130_fd_sc_hd__o21a_1 _10177_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_03521_),
    .B1(_03206_),
    .X(_03529_));
 sky130_fd_sc_hd__xor2_2 _10178_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__xnor2_2 _10179_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__o21ai_1 _10180_ (.A1(_03519_),
    .A2(_03526_),
    .B1(_03524_),
    .Y(_03532_));
 sky130_fd_sc_hd__nor2_1 _10181_ (.A(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__a21o_1 _10182_ (.A1(_03531_),
    .A2(_03532_),
    .B1(_03183_),
    .X(_03534_));
 sky130_fd_sc_hd__o221a_1 _10183_ (.A1(_03191_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_03533_),
    .B2(_03534_),
    .C1(_03258_),
    .X(_00412_));
 sky130_fd_sc_hd__clkbuf_4 _10184_ (.A(_01765_),
    .X(_03535_));
 sky130_fd_sc_hd__or3_4 _10185_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .C(_03521_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_1 _10186_ (.A(_03207_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__xor2_2 _10187_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03537_),
    .X(_03538_));
 sky130_fd_sc_hd__xnor2_2 _10188_ (.A(_03105_),
    .B(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__a22o_1 _10189_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_03523_),
    .B1(_03530_),
    .B2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_03540_));
 sky130_fd_sc_hd__o21ai_1 _10190_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_03530_),
    .B1(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__o31a_1 _10191_ (.A1(_03519_),
    .A2(_03526_),
    .A3(_03531_),
    .B1(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__xor2_1 _10192_ (.A(_03539_),
    .B(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _10193_ (.A0(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A1(_03543_),
    .S(_03185_),
    .X(_03544_));
 sky130_fd_sc_hd__and2_1 _10194_ (.A(_03535_),
    .B(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(_03545_),
    .X(_00413_));
 sky130_fd_sc_hd__o21a_1 _10196_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_03536_),
    .B1(_03206_),
    .X(_03546_));
 sky130_fd_sc_hd__xor2_2 _10197_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__xnor2_1 _10198_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__nor2_1 _10199_ (.A(_03105_),
    .B(_03538_),
    .Y(_03549_));
 sky130_fd_sc_hd__o21ba_1 _10200_ (.A1(_03539_),
    .A2(_03542_),
    .B1_N(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__xor2_1 _10201_ (.A(_03548_),
    .B(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__or2_1 _10202_ (.A(_03190_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(_03552_));
 sky130_fd_sc_hd__o211a_1 _10203_ (.A1(_03389_),
    .A2(_03551_),
    .B1(_03552_),
    .C1(_03515_),
    .X(_00414_));
 sky130_fd_sc_hd__a21o_1 _10204_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_03547_),
    .B1(_03549_),
    .X(_03553_));
 sky130_fd_sc_hd__o21ai_1 _10205_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_03547_),
    .B1(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__or4_1 _10206_ (.A(_03526_),
    .B(_03531_),
    .C(_03539_),
    .D(_03548_),
    .X(_03555_));
 sky130_fd_sc_hd__a21o_1 _10207_ (.A1(_03517_),
    .A2(_03518_),
    .B1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__or3_1 _10208_ (.A(_03539_),
    .B(_03541_),
    .C(_03548_),
    .X(_03557_));
 sky130_fd_sc_hd__inv_2 _10209_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .Y(_03558_));
 sky130_fd_sc_hd__o31a_1 _10210_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A3(_03536_),
    .B1(_03207_),
    .X(_03559_));
 sky130_fd_sc_hd__xnor2_1 _10211_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__or2_1 _10212_ (.A(_03558_),
    .B(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _10213_ (.A(_03558_),
    .B(_03560_),
    .Y(_03562_));
 sky130_fd_sc_hd__nand2_1 _10214_ (.A(_03561_),
    .B(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__a31o_1 _10215_ (.A1(_03554_),
    .A2(_03556_),
    .A3(_03557_),
    .B1(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__nand4_1 _10216_ (.A(_03563_),
    .B(_03554_),
    .C(_03556_),
    .D(_03557_),
    .Y(_03565_));
 sky130_fd_sc_hd__and2_1 _10217_ (.A(_03564_),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__or2_1 _10218_ (.A(_03190_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_03567_));
 sky130_fd_sc_hd__o211a_1 _10219_ (.A1(_03389_),
    .A2(_03566_),
    .B1(_03567_),
    .C1(_03515_),
    .X(_00415_));
 sky130_fd_sc_hd__clkbuf_4 _10220_ (.A(_01455_),
    .X(_03568_));
 sky130_fd_sc_hd__nor4_2 _10221_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .D(_03536_),
    .Y(_03569_));
 sky130_fd_sc_hd__nor2_1 _10222_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A1(_03570_),
    .S(_03207_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_4 _10224_ (.A(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__and2_1 _10225_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_03569_),
    .X(_03573_));
 sky130_fd_sc_hd__or3_2 _10226_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03572_),
    .C(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__inv_2 _10227_ (.A(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__o21ai_1 _10228_ (.A1(_03572_),
    .A2(_03573_),
    .B1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .Y(_03576_));
 sky130_fd_sc_hd__nand2_1 _10229_ (.A(_03561_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__or2b_1 _10230_ (.A(_03577_),
    .B_N(_03564_),
    .X(_03578_));
 sky130_fd_sc_hd__and2_1 _10231_ (.A(_03574_),
    .B(_03576_),
    .X(_03579_));
 sky130_fd_sc_hd__a21o_1 _10232_ (.A1(_03561_),
    .A2(_03564_),
    .B1(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__o211ai_1 _10233_ (.A1(_03575_),
    .A2(_03578_),
    .B1(_03580_),
    .C1(_03191_),
    .Y(_03581_));
 sky130_fd_sc_hd__o211a_1 _10234_ (.A1(_03189_),
    .A2(net437),
    .B1(_03568_),
    .C1(_03581_),
    .X(_00416_));
 sky130_fd_sc_hd__and2_1 _10235_ (.A(_03201_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_03582_));
 sky130_fd_sc_hd__xnor2_1 _10236_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_03572_),
    .Y(_03583_));
 sky130_fd_sc_hd__and3b_1 _10237_ (.A_N(_03583_),
    .B(_03578_),
    .C(_03574_),
    .X(_03584_));
 sky130_fd_sc_hd__a21bo_1 _10238_ (.A1(_03574_),
    .A2(_03578_),
    .B1_N(_03583_),
    .X(_03585_));
 sky130_fd_sc_hd__and3b_1 _10239_ (.A_N(_03584_),
    .B(_03585_),
    .C(_03186_),
    .X(_03586_));
 sky130_fd_sc_hd__o21a_1 _10240_ (.A1(_03582_),
    .A2(_03586_),
    .B1(_02132_),
    .X(_00417_));
 sky130_fd_sc_hd__a21o_1 _10241_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_03572_),
    .B1(_03584_),
    .X(_03587_));
 sky130_fd_sc_hd__xnor2_1 _10242_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_03572_),
    .Y(_03588_));
 sky130_fd_sc_hd__xnor2_1 _10243_ (.A(_03587_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__or2_1 _10244_ (.A(_03190_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(_03590_));
 sky130_fd_sc_hd__o211a_1 _10245_ (.A1(_03183_),
    .A2(_03589_),
    .B1(_03590_),
    .C1(_03515_),
    .X(_00418_));
 sky130_fd_sc_hd__and2_1 _10246_ (.A(_03201_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .X(_03591_));
 sky130_fd_sc_hd__nor2_1 _10247_ (.A(_03583_),
    .B(_03588_),
    .Y(_03592_));
 sky130_fd_sc_hd__and3b_1 _10248_ (.A_N(_03564_),
    .B(_03579_),
    .C(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__a32o_1 _10249_ (.A1(_03574_),
    .A2(_03577_),
    .A3(_03592_),
    .B1(_03572_),
    .B2(_03390_),
    .X(_03594_));
 sky130_fd_sc_hd__xor2_1 _10250_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03572_),
    .X(_03595_));
 sky130_fd_sc_hd__o21a_1 _10251_ (.A1(_03593_),
    .A2(_03594_),
    .B1(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__or3_1 _10252_ (.A(_03595_),
    .B(_03593_),
    .C(_03594_),
    .X(_03597_));
 sky130_fd_sc_hd__and3b_1 _10253_ (.A_N(_03596_),
    .B(_03597_),
    .C(_03186_),
    .X(_03598_));
 sky130_fd_sc_hd__o21a_1 _10254_ (.A1(_03591_),
    .A2(_03598_),
    .B1(_02132_),
    .X(_00419_));
 sky130_fd_sc_hd__a21o_1 _10255_ (.A1(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_03572_),
    .B1(_03596_),
    .X(_03599_));
 sky130_fd_sc_hd__xnor2_1 _10256_ (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_03572_),
    .Y(_03600_));
 sky130_fd_sc_hd__nor2_1 _10257_ (.A(_03599_),
    .B(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__a21o_1 _10258_ (.A1(_03599_),
    .A2(_03600_),
    .B1(_03201_),
    .X(_03602_));
 sky130_fd_sc_hd__o221a_1 _10259_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_03237_),
    .B1(_03601_),
    .B2(_03602_),
    .C1(_03258_),
    .X(_00420_));
 sky130_fd_sc_hd__and2_1 _10260_ (.A(_03186_),
    .B(_02310_),
    .X(_03603_));
 sky130_fd_sc_hd__clkbuf_1 _10261_ (.A(_03603_),
    .X(_00421_));
 sky130_fd_sc_hd__inv_2 _10262_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_03604_));
 sky130_fd_sc_hd__clkbuf_4 _10263_ (.A(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__clkbuf_4 _10264_ (.A(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__clkbuf_4 _10265_ (.A(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__buf_2 _10266_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03608_));
 sky130_fd_sc_hd__buf_2 _10267_ (.A(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__or2_1 _10268_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__o211a_1 _10269_ (.A1(_03607_),
    .A2(net216),
    .B1(_03568_),
    .C1(_03610_),
    .X(_00422_));
 sky130_fd_sc_hd__or2_1 _10270_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_03609_),
    .X(_03611_));
 sky130_fd_sc_hd__o211a_1 _10271_ (.A1(_03607_),
    .A2(net132),
    .B1(_03568_),
    .C1(_03611_),
    .X(_00423_));
 sky130_fd_sc_hd__or2_1 _10272_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B(_03609_),
    .X(_03612_));
 sky130_fd_sc_hd__o211a_1 _10273_ (.A1(_03607_),
    .A2(net141),
    .B1(_03568_),
    .C1(_03612_),
    .X(_00424_));
 sky130_fd_sc_hd__or2_1 _10274_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(_03609_),
    .X(_03613_));
 sky130_fd_sc_hd__o211a_1 _10275_ (.A1(_03607_),
    .A2(net136),
    .B1(_03568_),
    .C1(_03613_),
    .X(_00425_));
 sky130_fd_sc_hd__or2_1 _10276_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(_03609_),
    .X(_03614_));
 sky130_fd_sc_hd__o211a_1 _10277_ (.A1(_03607_),
    .A2(net130),
    .B1(_03568_),
    .C1(_03614_),
    .X(_00426_));
 sky130_fd_sc_hd__or2_1 _10278_ (.A(net265),
    .B(_03609_),
    .X(_03615_));
 sky130_fd_sc_hd__o211a_1 _10279_ (.A1(_03607_),
    .A2(net266),
    .B1(_03568_),
    .C1(_03615_),
    .X(_00427_));
 sky130_fd_sc_hd__or2_1 _10280_ (.A(net234),
    .B(_03609_),
    .X(_03616_));
 sky130_fd_sc_hd__o211a_1 _10281_ (.A1(_03607_),
    .A2(net254),
    .B1(_03568_),
    .C1(_03616_),
    .X(_00428_));
 sky130_fd_sc_hd__or2_1 _10282_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_03609_),
    .X(_03617_));
 sky130_fd_sc_hd__o211a_1 _10283_ (.A1(_03607_),
    .A2(net126),
    .B1(_03568_),
    .C1(_03617_),
    .X(_00429_));
 sky130_fd_sc_hd__or2_1 _10284_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_03609_),
    .X(_03618_));
 sky130_fd_sc_hd__o211a_1 _10285_ (.A1(_03607_),
    .A2(net124),
    .B1(_03568_),
    .C1(_03618_),
    .X(_00430_));
 sky130_fd_sc_hd__clkbuf_4 _10286_ (.A(_01251_),
    .X(_03619_));
 sky130_fd_sc_hd__clkbuf_4 _10287_ (.A(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_2 _10288_ (.A(_03608_),
    .X(_03621_));
 sky130_fd_sc_hd__or2_1 _10289_ (.A(net158),
    .B(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__o211a_1 _10290_ (.A1(_03607_),
    .A2(net298),
    .B1(_03620_),
    .C1(_03622_),
    .X(_00431_));
 sky130_fd_sc_hd__clkbuf_4 _10291_ (.A(_03606_),
    .X(_03623_));
 sky130_fd_sc_hd__or2_1 _10292_ (.A(_03609_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(_03624_));
 sky130_fd_sc_hd__o211a_1 _10293_ (.A1(_03623_),
    .A2(net252),
    .B1(_03620_),
    .C1(_03624_),
    .X(_00432_));
 sky130_fd_sc_hd__buf_2 _10294_ (.A(_03608_),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_4 _10295_ (.A(_03608_),
    .X(_03626_));
 sky130_fd_sc_hd__nand2_1 _10296_ (.A(_03626_),
    .B(net377),
    .Y(_03627_));
 sky130_fd_sc_hd__o211a_1 _10297_ (.A1(_03625_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_03620_),
    .C1(_03627_),
    .X(_00433_));
 sky130_fd_sc_hd__nand2_1 _10298_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_03628_));
 sky130_fd_sc_hd__or2_1 _10299_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(_03629_));
 sky130_fd_sc_hd__a21oi_2 _10300_ (.A1(_03628_),
    .A2(_03629_),
    .B1(_03280_),
    .Y(_03630_));
 sky130_fd_sc_hd__clkbuf_4 _10301_ (.A(_03605_),
    .X(_03631_));
 sky130_fd_sc_hd__a31o_1 _10302_ (.A1(_03280_),
    .A2(_03628_),
    .A3(_03629_),
    .B1(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_4 _10303_ (.A(_02308_),
    .X(_03633_));
 sky130_fd_sc_hd__o221a_1 _10304_ (.A1(_03625_),
    .A2(net592),
    .B1(_03630_),
    .B2(_03632_),
    .C1(_03633_),
    .X(_00434_));
 sky130_fd_sc_hd__and3_1 _10305_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(_03634_));
 sky130_fd_sc_hd__a21oi_1 _10306_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .Y(_03635_));
 sky130_fd_sc_hd__or2_1 _10307_ (.A(_03634_),
    .B(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__nor2_1 _10308_ (.A(_03630_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__a21o_1 _10309_ (.A1(_03630_),
    .A2(_03636_),
    .B1(_03606_),
    .X(_03638_));
 sky130_fd_sc_hd__o221a_1 _10310_ (.A1(_03625_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B1(_03637_),
    .B2(_03638_),
    .C1(_03633_),
    .X(_00435_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(_03280_),
    .B(_03634_),
    .Y(_03639_));
 sky130_fd_sc_hd__o31a_1 _10312_ (.A1(_03280_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(_03629_),
    .B1(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__and2_1 _10313_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_4 _10314_ (.A(_03608_),
    .X(_03642_));
 sky130_fd_sc_hd__o21ai_1 _10315_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_03640_),
    .B1(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__o221a_1 _10316_ (.A1(_03625_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_03641_),
    .B2(_03643_),
    .C1(_03633_),
    .X(_00436_));
 sky130_fd_sc_hd__or3_1 _10317_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_03629_),
    .X(_03644_));
 sky130_fd_sc_hd__nand2_1 _10318_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_03634_),
    .Y(_03645_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(_03644_),
    .A1(_03645_),
    .S(_03280_),
    .X(_03646_));
 sky130_fd_sc_hd__and2_1 _10320_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__o21ai_1 _10321_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_03646_),
    .B1(_03642_),
    .Y(_03648_));
 sky130_fd_sc_hd__o221a_1 _10322_ (.A1(_03625_),
    .A2(net501),
    .B1(_03647_),
    .B2(_03648_),
    .C1(_03633_),
    .X(_00437_));
 sky130_fd_sc_hd__inv_2 _10323_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_03649_));
 sky130_fd_sc_hd__buf_2 _10324_ (.A(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_4 _10325_ (.A(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__o21ai_1 _10326_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_03644_),
    .B1(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a31o_1 _10327_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A3(_03634_),
    .B1(_03651_),
    .X(_03653_));
 sky130_fd_sc_hd__inv_2 _10328_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .Y(_03654_));
 sky130_fd_sc_hd__a21oi_1 _10329_ (.A1(_03652_),
    .A2(_03653_),
    .B1(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__a31o_1 _10330_ (.A1(_03654_),
    .A2(_03652_),
    .A3(_03653_),
    .B1(_03631_),
    .X(_03656_));
 sky130_fd_sc_hd__o221a_1 _10331_ (.A1(_03625_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_03655_),
    .B2(_03656_),
    .C1(_03633_),
    .X(_00438_));
 sky130_fd_sc_hd__and4_1 _10332_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .D(_03634_),
    .X(_03657_));
 sky130_fd_sc_hd__or3_1 _10333_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_03644_),
    .X(_03658_));
 sky130_fd_sc_hd__inv_2 _10334_ (.A(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(_03657_),
    .A1(_03659_),
    .S(_03651_),
    .X(_03660_));
 sky130_fd_sc_hd__xnor2_1 _10336_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__nand2_1 _10337_ (.A(_03642_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__o211a_1 _10338_ (.A1(_03625_),
    .A2(net428),
    .B1(_03620_),
    .C1(_03662_),
    .X(_00439_));
 sky130_fd_sc_hd__o21a_1 _10339_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_03658_),
    .B1(_03651_),
    .X(_03663_));
 sky130_fd_sc_hd__a21o_1 _10340_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_03657_),
    .B1(_03651_),
    .X(_03664_));
 sky130_fd_sc_hd__or2b_1 _10341_ (.A(_03663_),
    .B_N(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__nor2_1 _10342_ (.A(net526),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__a21o_1 _10343_ (.A1(net537),
    .A2(_03665_),
    .B1(_03606_),
    .X(_03667_));
 sky130_fd_sc_hd__o221a_1 _10344_ (.A1(_03626_),
    .A2(net444),
    .B1(_03666_),
    .B2(_03667_),
    .C1(_03633_),
    .X(_00440_));
 sky130_fd_sc_hd__a21oi_1 _10345_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_03664_),
    .B1(_03663_),
    .Y(_03668_));
 sky130_fd_sc_hd__buf_2 _10346_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_03669_));
 sky130_fd_sc_hd__or2_1 _10347_ (.A(_03621_),
    .B(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__o211a_1 _10348_ (.A1(_03623_),
    .A2(_03668_),
    .B1(_03670_),
    .C1(_03515_),
    .X(_00441_));
 sky130_fd_sc_hd__inv_2 _10349_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .Y(_03671_));
 sky130_fd_sc_hd__nor2_1 _10350_ (.A(_03671_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_03672_));
 sky130_fd_sc_hd__a21o_1 _10351_ (.A1(_03671_),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_03606_),
    .X(_03673_));
 sky130_fd_sc_hd__o221a_1 _10352_ (.A1(_03626_),
    .A2(net569),
    .B1(_03672_),
    .B2(_03673_),
    .C1(_03633_),
    .X(_00442_));
 sky130_fd_sc_hd__and2b_1 _10353_ (.A_N(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_03674_));
 sky130_fd_sc_hd__xnor2_1 _10354_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__xnor2_1 _10355_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__xor2_1 _10356_ (.A(_03672_),
    .B(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__or2_1 _10357_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_03678_));
 sky130_fd_sc_hd__o211a_1 _10358_ (.A1(_03623_),
    .A2(_03677_),
    .B1(_03678_),
    .C1(_03515_),
    .X(_00443_));
 sky130_fd_sc_hd__and2_1 _10359_ (.A(_03631_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .X(_03679_));
 sky130_fd_sc_hd__inv_2 _10360_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_03680_));
 sky130_fd_sc_hd__a21oi_1 _10361_ (.A1(_03680_),
    .A2(_03671_),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_03681_));
 sky130_fd_sc_hd__xnor2_1 _10362_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__or2_1 _10363_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__nand2_1 _10364_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_03682_),
    .Y(_03684_));
 sky130_fd_sc_hd__and2_1 _10365_ (.A(_03683_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__nand2_1 _10366_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_03675_),
    .Y(_03686_));
 sky130_fd_sc_hd__o21ai_1 _10367_ (.A1(_03672_),
    .A2(_03676_),
    .B1(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__o21ai_1 _10368_ (.A1(_03685_),
    .A2(_03687_),
    .B1(_03642_),
    .Y(_03688_));
 sky130_fd_sc_hd__a21oi_1 _10369_ (.A1(_03685_),
    .A2(_03687_),
    .B1(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__o21a_1 _10370_ (.A1(_03679_),
    .A2(_03689_),
    .B1(_02132_),
    .X(_00444_));
 sky130_fd_sc_hd__o31a_1 _10371_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A3(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B1(_03650_),
    .X(_03690_));
 sky130_fd_sc_hd__xnor2_1 _10372_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__and2_1 _10373_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__nor2_1 _10374_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__nor2_1 _10375_ (.A(_03692_),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__a21bo_1 _10376_ (.A1(_03683_),
    .A2(_03687_),
    .B1_N(_03684_),
    .X(_03695_));
 sky130_fd_sc_hd__xor2_1 _10377_ (.A(_03694_),
    .B(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__mux2_1 _10378_ (.A0(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_03696_),
    .S(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03697_));
 sky130_fd_sc_hd__and2_1 _10379_ (.A(_03535_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _10380_ (.A(_03698_),
    .X(_00445_));
 sky130_fd_sc_hd__a21o_1 _10381_ (.A1(_03694_),
    .A2(_03695_),
    .B1(_03692_),
    .X(_03699_));
 sky130_fd_sc_hd__nor4_1 _10382_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .C(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .D(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_1 _10383_ (.A(_03280_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__xnor2_1 _10384_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__and2_1 _10385_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__nor2_1 _10386_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__or2_1 _10387_ (.A(_03703_),
    .B(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__xnor2_1 _10388_ (.A(_03699_),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__or2_1 _10389_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(_03707_));
 sky130_fd_sc_hd__o211a_1 _10390_ (.A1(_03623_),
    .A2(_03706_),
    .B1(_03707_),
    .C1(_03515_),
    .X(_00446_));
 sky130_fd_sc_hd__inv_2 _10391_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .Y(_03708_));
 sky130_fd_sc_hd__or4_1 _10392_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .C(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .D(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_03709_));
 sky130_fd_sc_hd__o21a_1 _10393_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_03709_),
    .B1(_03650_),
    .X(_03710_));
 sky130_fd_sc_hd__xnor2_1 _10394_ (.A(_03708_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__and2b_1 _10395_ (.A_N(_03711_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_03712_));
 sky130_fd_sc_hd__or2b_1 _10396_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B_N(_03711_),
    .X(_03713_));
 sky130_fd_sc_hd__or2b_1 _10397_ (.A(_03712_),
    .B_N(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__inv_2 _10398_ (.A(_03705_),
    .Y(_03715_));
 sky130_fd_sc_hd__a21o_1 _10399_ (.A1(_03699_),
    .A2(_03715_),
    .B1(_03703_),
    .X(_03716_));
 sky130_fd_sc_hd__and2_1 _10400_ (.A(_03714_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__o21ai_1 _10401_ (.A1(_03714_),
    .A2(_03716_),
    .B1(_03642_),
    .Y(_03718_));
 sky130_fd_sc_hd__o221a_1 _10402_ (.A1(_03626_),
    .A2(net393),
    .B1(_03717_),
    .B2(_03718_),
    .C1(_03633_),
    .X(_00447_));
 sky130_fd_sc_hd__nor2_1 _10403_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .Y(_03719_));
 sky130_fd_sc_hd__a21oi_1 _10404_ (.A1(net117),
    .A2(_03719_),
    .B1(_03280_),
    .Y(_03720_));
 sky130_fd_sc_hd__xnor2_1 _10405_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__and2_1 _10406_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__nor2_1 _10407_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03721_),
    .Y(_03723_));
 sky130_fd_sc_hd__nor2_2 _10408_ (.A(_03722_),
    .B(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__nor2_1 _10409_ (.A(_03705_),
    .B(_03714_),
    .Y(_03725_));
 sky130_fd_sc_hd__o21a_1 _10410_ (.A1(_03703_),
    .A2(_03712_),
    .B1(_03713_),
    .X(_03726_));
 sky130_fd_sc_hd__a21o_1 _10411_ (.A1(_03699_),
    .A2(_03725_),
    .B1(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__nand2_1 _10412_ (.A(_03724_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__o21a_1 _10413_ (.A1(_03724_),
    .A2(_03727_),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03729_));
 sky130_fd_sc_hd__a22o_1 _10414_ (.A1(_03605_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_03728_),
    .B2(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__and2_1 _10415_ (.A(_03535_),
    .B(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _10416_ (.A(_03731_),
    .X(_00448_));
 sky130_fd_sc_hd__a21oi_1 _10417_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_03650_),
    .B1(_03720_),
    .Y(_03732_));
 sky130_fd_sc_hd__xnor2_2 _10418_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__xnor2_2 _10419_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__a21oi_1 _10420_ (.A1(_03724_),
    .A2(_03727_),
    .B1(_03722_),
    .Y(_03735_));
 sky130_fd_sc_hd__xnor2_1 _10421_ (.A(_03734_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__or2_1 _10422_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_03737_));
 sky130_fd_sc_hd__o211a_1 _10423_ (.A1(_03623_),
    .A2(_03736_),
    .B1(_03737_),
    .C1(_03515_),
    .X(_00449_));
 sky130_fd_sc_hd__inv_2 _10424_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .Y(_03738_));
 sky130_fd_sc_hd__o21ba_1 _10425_ (.A1(_03738_),
    .A2(_03733_),
    .B1_N(_03722_),
    .X(_03739_));
 sky130_fd_sc_hd__a21oi_1 _10426_ (.A1(_03738_),
    .A2(_03733_),
    .B1(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__a31oi_2 _10427_ (.A1(_03724_),
    .A2(_03726_),
    .A3(_03734_),
    .B1(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand4_2 _10428_ (.A(_03699_),
    .B(_03724_),
    .C(_03725_),
    .D(_03734_),
    .Y(_03742_));
 sky130_fd_sc_hd__and2_1 _10429_ (.A(_03741_),
    .B(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__nor2_1 _10430_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .Y(_03744_));
 sky130_fd_sc_hd__a31o_1 _10431_ (.A1(net117),
    .A2(_03719_),
    .A3(_03744_),
    .B1(_03280_),
    .X(_03745_));
 sky130_fd_sc_hd__xor2_1 _10432_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _10433_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__or2_1 _10434_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03746_),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_1 _10435_ (.A(_03747_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__xor2_1 _10436_ (.A(_03743_),
    .B(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__or2_1 _10437_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_03751_));
 sky130_fd_sc_hd__o211a_1 _10438_ (.A1(_03623_),
    .A2(_03750_),
    .B1(_03751_),
    .C1(_03515_),
    .X(_00450_));
 sky130_fd_sc_hd__inv_2 _10439_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .Y(_03752_));
 sky130_fd_sc_hd__a21boi_1 _10440_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_03651_),
    .B1_N(_03745_),
    .Y(_03753_));
 sky130_fd_sc_hd__xnor2_2 _10441_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__xnor2_1 _10442_ (.A(_03752_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__o21ai_1 _10443_ (.A1(_03743_),
    .A2(_03749_),
    .B1(_03747_),
    .Y(_03756_));
 sky130_fd_sc_hd__nor2_1 _10444_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__a21o_1 _10445_ (.A1(_03755_),
    .A2(_03756_),
    .B1(_03631_),
    .X(_03758_));
 sky130_fd_sc_hd__o221a_1 _10446_ (.A1(_03626_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_03757_),
    .B2(_03758_),
    .C1(_03633_),
    .X(_00451_));
 sky130_fd_sc_hd__nor2_1 _10447_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .Y(_03759_));
 sky130_fd_sc_hd__and4_1 _10448_ (.A(net117),
    .B(_03719_),
    .C(_03744_),
    .D(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__nor2_1 _10449_ (.A(_03280_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__xnor2_1 _10450_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__or2_1 _10452_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03762_),
    .X(_03764_));
 sky130_fd_sc_hd__and2_1 _10453_ (.A(_03763_),
    .B(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__or2_1 _10454_ (.A(_03749_),
    .B(_03755_),
    .X(_03766_));
 sky130_fd_sc_hd__o21a_1 _10455_ (.A1(_03752_),
    .A2(_03754_),
    .B1(_03747_),
    .X(_03767_));
 sky130_fd_sc_hd__a21o_1 _10456_ (.A1(_03752_),
    .A2(_03754_),
    .B1(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__o21ai_1 _10457_ (.A1(_03743_),
    .A2(_03766_),
    .B1(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__xor2_1 _10458_ (.A(_03765_),
    .B(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A1(_03770_),
    .S(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03771_));
 sky130_fd_sc_hd__and2_1 _10460_ (.A(_03535_),
    .B(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_03772_),
    .X(_00452_));
 sky130_fd_sc_hd__or2b_1 _10462_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B_N(_03760_),
    .X(_03773_));
 sky130_fd_sc_hd__nand2_1 _10463_ (.A(_03651_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__xor2_2 _10464_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__xor2_1 _10465_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__a21bo_1 _10466_ (.A1(_03765_),
    .A2(_03769_),
    .B1_N(_03763_),
    .X(_03777_));
 sky130_fd_sc_hd__xor2_1 _10467_ (.A(_03776_),
    .B(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__or2_1 _10468_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_03779_));
 sky130_fd_sc_hd__clkbuf_4 _10469_ (.A(_01474_),
    .X(_03780_));
 sky130_fd_sc_hd__o211a_1 _10470_ (.A1(_03623_),
    .A2(_03778_),
    .B1(_03779_),
    .C1(_03780_),
    .X(_00453_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(_03765_),
    .B(_03776_),
    .Y(_03781_));
 sky130_fd_sc_hd__a211o_1 _10472_ (.A1(_03741_),
    .A2(_03742_),
    .B1(_03766_),
    .C1(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__a21bo_1 _10473_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_03775_),
    .B1_N(_03763_),
    .X(_03783_));
 sky130_fd_sc_hd__o21ai_2 _10474_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_03775_),
    .B1(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__or2_1 _10475_ (.A(_03768_),
    .B(_03781_),
    .X(_03785_));
 sky130_fd_sc_hd__o21ai_1 _10476_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_03773_),
    .B1(_03651_),
    .Y(_03786_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(_03786_),
    .A1(_03651_),
    .S(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_03787_));
 sky130_fd_sc_hd__or3b_1 _10478_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03773_),
    .C_N(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_03788_));
 sky130_fd_sc_hd__and3_1 _10479_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_03787_),
    .C(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__a21oi_1 _10480_ (.A1(_03787_),
    .A2(_03788_),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .Y(_03790_));
 sky130_fd_sc_hd__or2_1 _10481_ (.A(_03789_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__a31oi_4 _10482_ (.A1(_03782_),
    .A2(_03784_),
    .A3(_03785_),
    .B1(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__and4_1 _10483_ (.A(_03791_),
    .B(_03782_),
    .C(_03784_),
    .D(_03785_),
    .X(_03793_));
 sky130_fd_sc_hd__nor2_1 _10484_ (.A(_03792_),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__or2_1 _10485_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_03795_));
 sky130_fd_sc_hd__o211a_1 _10486_ (.A1(_03623_),
    .A2(_03794_),
    .B1(_03795_),
    .C1(_03780_),
    .X(_00454_));
 sky130_fd_sc_hd__clkbuf_4 _10487_ (.A(_03787_),
    .X(_03796_));
 sky130_fd_sc_hd__xor2_1 _10488_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__o21ba_1 _10489_ (.A1(_03789_),
    .A2(_03792_),
    .B1_N(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__or3b_1 _10490_ (.A(_03789_),
    .B(_03792_),
    .C_N(_03797_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_1 _10491_ (.A(_03642_),
    .B(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__o221a_1 _10492_ (.A1(_03626_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_03798_),
    .B2(_03800_),
    .C1(_03633_),
    .X(_00455_));
 sky130_fd_sc_hd__inv_2 _10493_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .Y(_03801_));
 sky130_fd_sc_hd__nor2_1 _10494_ (.A(_03642_),
    .B(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__o21ai_1 _10495_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_03796_),
    .B1(_03792_),
    .Y(_03803_));
 sky130_fd_sc_hd__a21oi_1 _10496_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_03796_),
    .B1(_03789_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _10497_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03796_),
    .Y(_03805_));
 sky130_fd_sc_hd__or2_1 _10498_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03796_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_1 _10499_ (.A(_03805_),
    .B(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__a21bo_1 _10500_ (.A1(_03803_),
    .A2(_03804_),
    .B1_N(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__nand3b_1 _10501_ (.A_N(_03807_),
    .B(_03803_),
    .C(_03804_),
    .Y(_03809_));
 sky130_fd_sc_hd__and3_1 _10502_ (.A(_03642_),
    .B(_03808_),
    .C(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__o21a_1 _10503_ (.A1(_03802_),
    .A2(_03810_),
    .B1(_02132_),
    .X(_00456_));
 sky130_fd_sc_hd__xor2_1 _10504_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_03796_),
    .X(_03811_));
 sky130_fd_sc_hd__a21oi_1 _10505_ (.A1(_03805_),
    .A2(_03808_),
    .B1(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__a31o_1 _10506_ (.A1(_03805_),
    .A2(_03808_),
    .A3(_03811_),
    .B1(_03631_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_4 _10507_ (.A(_02308_),
    .X(_03814_));
 sky130_fd_sc_hd__o221a_1 _10508_ (.A1(_03626_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B1(_03812_),
    .B2(_03813_),
    .C1(_03814_),
    .X(_00457_));
 sky130_fd_sc_hd__or2_1 _10509_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03796_),
    .X(_03815_));
 sky130_fd_sc_hd__nand2_1 _10510_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03796_),
    .Y(_03816_));
 sky130_fd_sc_hd__and2_1 _10511_ (.A(_03815_),
    .B(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__and4_1 _10512_ (.A(_03792_),
    .B(_03797_),
    .C(_03807_),
    .D(_03811_),
    .X(_03818_));
 sky130_fd_sc_hd__o21a_1 _10513_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_03796_),
    .X(_03819_));
 sky130_fd_sc_hd__or3b_1 _10514_ (.A(_03818_),
    .B(_03819_),
    .C_N(_03804_),
    .X(_03820_));
 sky130_fd_sc_hd__nand2_1 _10515_ (.A(_03817_),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__o21a_1 _10516_ (.A1(_03817_),
    .A2(_03820_),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03822_));
 sky130_fd_sc_hd__a22o_1 _10517_ (.A1(_03605_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B1(_03821_),
    .B2(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_1 _10518_ (.A(_03535_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(_03824_),
    .X(_00458_));
 sky130_fd_sc_hd__xor2_1 _10520_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_03796_),
    .X(_03825_));
 sky130_fd_sc_hd__a21oi_1 _10521_ (.A1(_03816_),
    .A2(_03821_),
    .B1(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__a31o_1 _10522_ (.A1(_03816_),
    .A2(_03821_),
    .A3(_03825_),
    .B1(_03631_),
    .X(_03827_));
 sky130_fd_sc_hd__o221a_1 _10523_ (.A1(_03626_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B1(_03826_),
    .B2(_03827_),
    .C1(_03814_),
    .X(_00459_));
 sky130_fd_sc_hd__and2_1 _10524_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_03828_));
 sky130_fd_sc_hd__nor2_1 _10525_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .Y(_03829_));
 sky130_fd_sc_hd__o21ai_2 _10526_ (.A1(_03828_),
    .A2(_03829_),
    .B1(_03642_),
    .Y(_03830_));
 sky130_fd_sc_hd__o211a_1 _10527_ (.A1(_03625_),
    .A2(net455),
    .B1(_03620_),
    .C1(_03830_),
    .X(_00460_));
 sky130_fd_sc_hd__and2b_1 _10528_ (.A_N(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_03831_));
 sky130_fd_sc_hd__xnor2_1 _10529_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__xnor2_1 _10530_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__xor2_1 _10531_ (.A(_03828_),
    .B(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__or2_1 _10532_ (.A(_03621_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_03835_));
 sky130_fd_sc_hd__o211a_1 _10533_ (.A1(_03623_),
    .A2(_03834_),
    .B1(_03835_),
    .C1(_03780_),
    .X(_00461_));
 sky130_fd_sc_hd__inv_2 _10534_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_03836_));
 sky130_fd_sc_hd__o21a_1 _10535_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B1(_03649_),
    .X(_03837_));
 sky130_fd_sc_hd__xnor2_1 _10536_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__and2_1 _10537_ (.A(_03836_),
    .B(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__nor2_1 _10538_ (.A(_03836_),
    .B(_03838_),
    .Y(_03840_));
 sky130_fd_sc_hd__nor2_1 _10539_ (.A(_03839_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__and2b_1 _10540_ (.A_N(_03832_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_03842_));
 sky130_fd_sc_hd__a21o_1 _10541_ (.A1(_03828_),
    .A2(_03833_),
    .B1(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_03841_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__o21a_1 _10543_ (.A1(_03841_),
    .A2(_03843_),
    .B1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03845_));
 sky130_fd_sc_hd__a22o_1 _10544_ (.A1(_03605_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_03844_),
    .B2(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__and2_1 _10545_ (.A(_03535_),
    .B(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_1 _10546_ (.A(_03847_),
    .X(_00462_));
 sky130_fd_sc_hd__inv_2 _10547_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_03848_));
 sky130_fd_sc_hd__o31a_1 _10548_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A3(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B1(_03649_),
    .X(_03849_));
 sky130_fd_sc_hd__xnor2_1 _10549_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _10550_ (.A(_03848_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__inv_2 _10551_ (.A(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _10552_ (.A(_03836_),
    .B(_03838_),
    .Y(_03853_));
 sky130_fd_sc_hd__a21o_1 _10553_ (.A1(_03853_),
    .A2(_03843_),
    .B1(_03840_),
    .X(_03854_));
 sky130_fd_sc_hd__a21o_1 _10554_ (.A1(_03852_),
    .A2(_03854_),
    .B1(_03605_),
    .X(_03855_));
 sky130_fd_sc_hd__nor2_1 _10555_ (.A(_03852_),
    .B(_03854_),
    .Y(_03856_));
 sky130_fd_sc_hd__a2bb2o_1 _10556_ (.A1_N(_03855_),
    .A2_N(_03856_),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B2(_03605_),
    .X(_03857_));
 sky130_fd_sc_hd__and2_1 _10557_ (.A(_03535_),
    .B(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_1 _10558_ (.A(_03858_),
    .X(_00463_));
 sky130_fd_sc_hd__nor2_1 _10559_ (.A(_03848_),
    .B(_03850_),
    .Y(_03859_));
 sky130_fd_sc_hd__a21oi_2 _10560_ (.A1(_03852_),
    .A2(_03854_),
    .B1(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__inv_2 _10561_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_03861_));
 sky130_fd_sc_hd__or4_4 _10562_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .C(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .D(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_03862_));
 sky130_fd_sc_hd__nand2_1 _10563_ (.A(_03650_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__xnor2_1 _10564_ (.A(_03752_),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__or2_1 _10565_ (.A(_03861_),
    .B(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__nand2_1 _10566_ (.A(_03861_),
    .B(_03864_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _10567_ (.A(_03865_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__xor2_1 _10568_ (.A(_03860_),
    .B(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__or2_1 _10569_ (.A(_03621_),
    .B(net510),
    .X(_03869_));
 sky130_fd_sc_hd__o211a_1 _10570_ (.A1(_03623_),
    .A2(_03868_),
    .B1(_03869_),
    .C1(_03780_),
    .X(_00464_));
 sky130_fd_sc_hd__o21a_1 _10571_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_03862_),
    .B1(_03649_),
    .X(_03870_));
 sky130_fd_sc_hd__xor2_2 _10572_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__nand2_2 _10573_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__or2_1 _10574_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03871_),
    .X(_03873_));
 sky130_fd_sc_hd__o21a_1 _10575_ (.A1(_03860_),
    .A2(_03867_),
    .B1(_03865_),
    .X(_03874_));
 sky130_fd_sc_hd__a21oi_1 _10576_ (.A1(_03872_),
    .A2(_03873_),
    .B1(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__a31o_1 _10577_ (.A1(_03872_),
    .A2(_03873_),
    .A3(_03874_),
    .B1(_03631_),
    .X(_03876_));
 sky130_fd_sc_hd__o221a_1 _10578_ (.A1(_03626_),
    .A2(net405),
    .B1(_03875_),
    .B2(_03876_),
    .C1(_03814_),
    .X(_00465_));
 sky130_fd_sc_hd__nor2_1 _10579_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_03871_),
    .Y(_03877_));
 sky130_fd_sc_hd__or2_1 _10580_ (.A(_03877_),
    .B(_03874_),
    .X(_03878_));
 sky130_fd_sc_hd__or2_1 _10581_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_03879_));
 sky130_fd_sc_hd__o21a_1 _10582_ (.A1(_03862_),
    .A2(_03879_),
    .B1(_03649_),
    .X(_03880_));
 sky130_fd_sc_hd__xnor2_1 _10583_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__nor2_1 _10584_ (.A(_03680_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__and2_1 _10585_ (.A(_03680_),
    .B(_03881_),
    .X(_03883_));
 sky130_fd_sc_hd__or2_1 _10586_ (.A(_03882_),
    .B(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__a21o_1 _10587_ (.A1(_03872_),
    .A2(_03878_),
    .B1(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__a31oi_1 _10588_ (.A1(_03872_),
    .A2(_03878_),
    .A3(_03884_),
    .B1(_03605_),
    .Y(_03886_));
 sky130_fd_sc_hd__a22o_1 _10589_ (.A1(_03605_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1(_03885_),
    .B2(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__and2_1 _10590_ (.A(_03535_),
    .B(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_03888_),
    .X(_00466_));
 sky130_fd_sc_hd__a21o_1 _10592_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_03650_),
    .B1(_03880_),
    .X(_03889_));
 sky130_fd_sc_hd__xor2_1 _10593_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__and2_1 _10594_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__nor2_1 _10595_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_03890_),
    .Y(_03892_));
 sky130_fd_sc_hd__or2_1 _10596_ (.A(_03891_),
    .B(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__and2b_1 _10597_ (.A_N(_03882_),
    .B(_03885_),
    .X(_03894_));
 sky130_fd_sc_hd__xor2_1 _10598_ (.A(_03893_),
    .B(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__or2_1 _10599_ (.A(_03608_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_03896_));
 sky130_fd_sc_hd__o211a_1 _10600_ (.A1(_03606_),
    .A2(_03895_),
    .B1(_03896_),
    .C1(_03780_),
    .X(_00467_));
 sky130_fd_sc_hd__a21o_1 _10601_ (.A1(_03865_),
    .A2(_03872_),
    .B1(_03877_),
    .X(_03897_));
 sky130_fd_sc_hd__nor2_1 _10602_ (.A(_03882_),
    .B(_03891_),
    .Y(_03898_));
 sky130_fd_sc_hd__o32a_1 _10603_ (.A1(_03884_),
    .A2(_03897_),
    .A3(_03893_),
    .B1(_03898_),
    .B2(_03892_),
    .X(_03899_));
 sky130_fd_sc_hd__nand2_1 _10604_ (.A(_03872_),
    .B(_03873_),
    .Y(_03900_));
 sky130_fd_sc_hd__or2_1 _10605_ (.A(_03867_),
    .B(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__or4_1 _10606_ (.A(_03860_),
    .B(_03884_),
    .C(_03901_),
    .D(_03893_),
    .X(_03902_));
 sky130_fd_sc_hd__and2_1 _10607_ (.A(_03899_),
    .B(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__or2_1 _10608_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_03904_));
 sky130_fd_sc_hd__or3_1 _10609_ (.A(_03862_),
    .B(_03879_),
    .C(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__nand2_1 _10610_ (.A(_03650_),
    .B(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__xnor2_1 _10611_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_1 _10612_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__or2_1 _10613_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_03907_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _10614_ (.A(_03908_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__xor2_1 _10615_ (.A(_03903_),
    .B(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__or2_1 _10616_ (.A(_03608_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_03912_));
 sky130_fd_sc_hd__o211a_1 _10617_ (.A1(_03606_),
    .A2(_03911_),
    .B1(_03912_),
    .C1(_03780_),
    .X(_00468_));
 sky130_fd_sc_hd__o21a_1 _10618_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_03905_),
    .B1(_03650_),
    .X(_03913_));
 sky130_fd_sc_hd__xor2_2 _10619_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__xnor2_2 _10620_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__o21ai_1 _10621_ (.A1(_03903_),
    .A2(_03910_),
    .B1(_03908_),
    .Y(_03916_));
 sky130_fd_sc_hd__nor2_1 _10622_ (.A(_03915_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__a21o_1 _10623_ (.A1(_03915_),
    .A2(_03916_),
    .B1(_03631_),
    .X(_03918_));
 sky130_fd_sc_hd__o221a_1 _10624_ (.A1(_03626_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_03917_),
    .B2(_03918_),
    .C1(_03814_),
    .X(_00469_));
 sky130_fd_sc_hd__or2_1 _10625_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_03919_));
 sky130_fd_sc_hd__or4_4 _10626_ (.A(_03862_),
    .B(_03879_),
    .C(_03904_),
    .D(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__nand2_1 _10627_ (.A(_03650_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__xor2_1 _10628_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__nor2_1 _10629_ (.A(_03708_),
    .B(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__and2_1 _10630_ (.A(_03708_),
    .B(_03922_),
    .X(_03924_));
 sky130_fd_sc_hd__or2_1 _10631_ (.A(_03923_),
    .B(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__a22o_1 _10632_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_03907_),
    .B1(_03914_),
    .B2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_03926_));
 sky130_fd_sc_hd__o21ai_2 _10633_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_03914_),
    .B1(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__or3_1 _10634_ (.A(_03903_),
    .B(_03910_),
    .C(_03915_),
    .X(_03928_));
 sky130_fd_sc_hd__a31o_1 _10635_ (.A1(_03925_),
    .A2(_03927_),
    .A3(_03928_),
    .B1(_03604_),
    .X(_03929_));
 sky130_fd_sc_hd__a21oi_1 _10636_ (.A1(_03927_),
    .A2(_03928_),
    .B1(_03925_),
    .Y(_03930_));
 sky130_fd_sc_hd__a2bb2o_1 _10637_ (.A1_N(_03929_),
    .A2_N(_03930_),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B2(_03605_),
    .X(_03931_));
 sky130_fd_sc_hd__and2_1 _10638_ (.A(_03535_),
    .B(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_03932_),
    .X(_00470_));
 sky130_fd_sc_hd__o21a_1 _10640_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_03920_),
    .B1(_03650_),
    .X(_03933_));
 sky130_fd_sc_hd__xor2_1 _10641_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__and2_1 _10642_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__nor2_1 _10643_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__or2_1 _10644_ (.A(_03935_),
    .B(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__or2_1 _10645_ (.A(_03923_),
    .B(_03930_),
    .X(_03938_));
 sky130_fd_sc_hd__xnor2_1 _10646_ (.A(_03937_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__or2_1 _10647_ (.A(_03608_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(_03940_));
 sky130_fd_sc_hd__o211a_1 _10648_ (.A1(_03606_),
    .A2(_03939_),
    .B1(_03940_),
    .C1(_03780_),
    .X(_00471_));
 sky130_fd_sc_hd__nor3_1 _10649_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(_03920_),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2_1 _10650_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A1(_03942_),
    .S(_03651_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_2 _10652_ (.A(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__a21oi_1 _10653_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A2(_03941_),
    .B1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__xnor2_1 _10654_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__or4_1 _10655_ (.A(_03910_),
    .B(_03915_),
    .C(_03925_),
    .D(_03937_),
    .X(_03947_));
 sky130_fd_sc_hd__a21o_1 _10656_ (.A1(_03899_),
    .A2(_03902_),
    .B1(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__a21oi_1 _10657_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_03934_),
    .B1(_03923_),
    .Y(_03949_));
 sky130_fd_sc_hd__o32a_1 _10658_ (.A1(_03925_),
    .A2(_03927_),
    .A3(_03937_),
    .B1(_03949_),
    .B2(_03936_),
    .X(_03950_));
 sky130_fd_sc_hd__and2_1 _10659_ (.A(_03948_),
    .B(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__xnor2_1 _10660_ (.A(_03946_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__or2_1 _10661_ (.A(_03608_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_03953_));
 sky130_fd_sc_hd__o211a_1 _10662_ (.A1(_03606_),
    .A2(_03952_),
    .B1(_03953_),
    .C1(_03780_),
    .X(_00472_));
 sky130_fd_sc_hd__or2_1 _10663_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03944_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_1 _10664_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03944_),
    .Y(_03955_));
 sky130_fd_sc_hd__nand2_1 _10665_ (.A(_03954_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__and2b_1 _10666_ (.A_N(_03945_),
    .B(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_03957_));
 sky130_fd_sc_hd__a21bo_1 _10667_ (.A1(_03948_),
    .A2(_03950_),
    .B1_N(_03946_),
    .X(_03958_));
 sky130_fd_sc_hd__or2b_1 _10668_ (.A(_03957_),
    .B_N(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_03944_),
    .Y(_03960_));
 sky130_fd_sc_hd__and2b_1 _10670_ (.A_N(_03957_),
    .B(_03955_),
    .X(_03961_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_03958_),
    .B(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__nor2_1 _10672_ (.A(_03960_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__a211o_1 _10673_ (.A1(_03956_),
    .A2(_03959_),
    .B1(_03631_),
    .C1(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__o211a_1 _10674_ (.A1(_03625_),
    .A2(net408),
    .B1(_03620_),
    .C1(_03964_),
    .X(_00473_));
 sky130_fd_sc_hd__nand2_1 _10675_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_03944_),
    .Y(_03965_));
 sky130_fd_sc_hd__or2_1 _10676_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_03943_),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _10677_ (.A(_03965_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__nand2_1 _10678_ (.A(_03954_),
    .B(_03962_),
    .Y(_03968_));
 sky130_fd_sc_hd__xor2_1 _10679_ (.A(_03967_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A1(_03969_),
    .S(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03970_));
 sky130_fd_sc_hd__and2_1 _10681_ (.A(_03535_),
    .B(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__clkbuf_1 _10682_ (.A(_03971_),
    .X(_00474_));
 sky130_fd_sc_hd__xnor2_1 _10683_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_03944_),
    .Y(_03972_));
 sky130_fd_sc_hd__o21ai_1 _10684_ (.A1(_03967_),
    .A2(_03968_),
    .B1(_03965_),
    .Y(_03973_));
 sky130_fd_sc_hd__xnor2_1 _10685_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__or2_1 _10686_ (.A(_03608_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(_03975_));
 sky130_fd_sc_hd__o211a_1 _10687_ (.A1(_03606_),
    .A2(_03974_),
    .B1(_03975_),
    .C1(_03780_),
    .X(_00475_));
 sky130_fd_sc_hd__clkbuf_4 _10688_ (.A(_01765_),
    .X(_03976_));
 sky130_fd_sc_hd__or2_1 _10689_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03944_),
    .X(_03977_));
 sky130_fd_sc_hd__nand2_1 _10690_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_03944_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _10691_ (.A(_03977_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__or2_1 _10692_ (.A(_03967_),
    .B(_03972_),
    .X(_03980_));
 sky130_fd_sc_hd__or3_1 _10693_ (.A(_03958_),
    .B(_03956_),
    .C(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__or3_1 _10694_ (.A(_03960_),
    .B(_03961_),
    .C(_03980_),
    .X(_03982_));
 sky130_fd_sc_hd__o21ai_1 _10695_ (.A1(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_03944_),
    .Y(_03983_));
 sky130_fd_sc_hd__and3_1 _10696_ (.A(_03981_),
    .B(_03982_),
    .C(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__xor2_1 _10697_ (.A(_03979_),
    .B(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A1(_03985_),
    .S(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03986_));
 sky130_fd_sc_hd__and2_1 _10699_ (.A(_03976_),
    .B(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_03987_),
    .X(_00476_));
 sky130_fd_sc_hd__or2_1 _10701_ (.A(_03979_),
    .B(_03984_),
    .X(_03988_));
 sky130_fd_sc_hd__xor2_1 _10702_ (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_03944_),
    .X(_03989_));
 sky130_fd_sc_hd__a21oi_1 _10703_ (.A1(_03978_),
    .A2(_03988_),
    .B1(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__a31o_1 _10704_ (.A1(_03978_),
    .A2(_03988_),
    .A3(_03989_),
    .B1(_03631_),
    .X(_03991_));
 sky130_fd_sc_hd__o221a_1 _10705_ (.A1(net535),
    .A2(_03625_),
    .B1(_03990_),
    .B2(_03991_),
    .C1(_03814_),
    .X(_00477_));
 sky130_fd_sc_hd__and2_1 _10706_ (.A(_03642_),
    .B(_02310_),
    .X(_03992_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(_03992_),
    .X(_00478_));
 sky130_fd_sc_hd__inv_2 _10708_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_03993_));
 sky130_fd_sc_hd__clkbuf_4 _10709_ (.A(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_4 _10710_ (.A(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__buf_4 _10711_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_4 _10712_ (.A(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__or2_1 _10713_ (.A(net157),
    .B(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__o211a_1 _10714_ (.A1(_03995_),
    .A2(net283),
    .B1(_03620_),
    .C1(_03998_),
    .X(_00479_));
 sky130_fd_sc_hd__buf_2 _10715_ (.A(_03996_),
    .X(_03999_));
 sky130_fd_sc_hd__or2_1 _10716_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__o211a_1 _10717_ (.A1(_03995_),
    .A2(net240),
    .B1(_03620_),
    .C1(_04000_),
    .X(_00480_));
 sky130_fd_sc_hd__or2_1 _10718_ (.A(net223),
    .B(_03999_),
    .X(_04001_));
 sky130_fd_sc_hd__o211a_1 _10719_ (.A1(_03995_),
    .A2(net225),
    .B1(_03620_),
    .C1(_04001_),
    .X(_00481_));
 sky130_fd_sc_hd__or2_1 _10720_ (.A(net175),
    .B(_03999_),
    .X(_04002_));
 sky130_fd_sc_hd__o211a_1 _10721_ (.A1(_03995_),
    .A2(net277),
    .B1(_03620_),
    .C1(_04002_),
    .X(_00482_));
 sky130_fd_sc_hd__clkbuf_4 _10722_ (.A(_03619_),
    .X(_04003_));
 sky130_fd_sc_hd__or2_1 _10723_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(_03999_),
    .X(_04004_));
 sky130_fd_sc_hd__o211a_1 _10724_ (.A1(_03995_),
    .A2(net186),
    .B1(_04003_),
    .C1(_04004_),
    .X(_00483_));
 sky130_fd_sc_hd__or2_1 _10725_ (.A(net261),
    .B(_03999_),
    .X(_04005_));
 sky130_fd_sc_hd__o211a_1 _10726_ (.A1(_03995_),
    .A2(net265),
    .B1(_04003_),
    .C1(_04005_),
    .X(_00484_));
 sky130_fd_sc_hd__or2_1 _10727_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_03999_),
    .X(_04006_));
 sky130_fd_sc_hd__o211a_1 _10728_ (.A1(_03995_),
    .A2(net234),
    .B1(_04003_),
    .C1(_04006_),
    .X(_00485_));
 sky130_fd_sc_hd__or2_1 _10729_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_03999_),
    .X(_04007_));
 sky130_fd_sc_hd__o211a_1 _10730_ (.A1(_03995_),
    .A2(net179),
    .B1(_04003_),
    .C1(_04007_),
    .X(_00486_));
 sky130_fd_sc_hd__or2_1 _10731_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_03999_),
    .X(_04008_));
 sky130_fd_sc_hd__o211a_1 _10732_ (.A1(_03995_),
    .A2(net172),
    .B1(_04003_),
    .C1(_04008_),
    .X(_00487_));
 sky130_fd_sc_hd__or2_1 _10733_ (.A(_03997_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(_04009_));
 sky130_fd_sc_hd__o211a_1 _10734_ (.A1(_03995_),
    .A2(net158),
    .B1(_04003_),
    .C1(_04009_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_2 _10735_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_4 _10736_ (.A(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__clkbuf_4 _10737_ (.A(_04010_),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_1 _10738_ (.A(_04012_),
    .B(net258),
    .Y(_04013_));
 sky130_fd_sc_hd__o211a_1 _10739_ (.A1(_04011_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B1(_04003_),
    .C1(_04013_),
    .X(_00489_));
 sky130_fd_sc_hd__nand2_1 _10740_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .Y(_04014_));
 sky130_fd_sc_hd__or2_1 _10741_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(_04015_));
 sky130_fd_sc_hd__a21oi_1 _10742_ (.A1(_04014_),
    .A2(_04015_),
    .B1(_03669_),
    .Y(_04016_));
 sky130_fd_sc_hd__a31o_1 _10743_ (.A1(_03669_),
    .A2(_04014_),
    .A3(_04015_),
    .B1(_03994_),
    .X(_04017_));
 sky130_fd_sc_hd__o221a_1 _10744_ (.A1(_04011_),
    .A2(net562),
    .B1(_04016_),
    .B2(_04017_),
    .C1(_03814_),
    .X(_00490_));
 sky130_fd_sc_hd__and3_1 _10745_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(_04018_));
 sky130_fd_sc_hd__a21oi_1 _10746_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .Y(_04019_));
 sky130_fd_sc_hd__or2_1 _10747_ (.A(_04018_),
    .B(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__nor2_1 _10748_ (.A(_04016_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21o_1 _10749_ (.A1(_04016_),
    .A2(_04020_),
    .B1(_03994_),
    .X(_04022_));
 sky130_fd_sc_hd__o221a_1 _10750_ (.A1(_04011_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_04021_),
    .B2(_04022_),
    .C1(_03814_),
    .X(_00491_));
 sky130_fd_sc_hd__clkbuf_4 _10751_ (.A(_04010_),
    .X(_04023_));
 sky130_fd_sc_hd__nand2_1 _10752_ (.A(_03669_),
    .B(_04018_),
    .Y(_04024_));
 sky130_fd_sc_hd__o31a_1 _10753_ (.A1(_03669_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A3(_04015_),
    .B1(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__and2_1 _10754_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__o21ai_1 _10755_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_04025_),
    .B1(_04012_),
    .Y(_04027_));
 sky130_fd_sc_hd__o221a_1 _10756_ (.A1(_04023_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B1(_04026_),
    .B2(_04027_),
    .C1(_03814_),
    .X(_00492_));
 sky130_fd_sc_hd__or3_1 _10757_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_04015_),
    .X(_04028_));
 sky130_fd_sc_hd__nand2_1 _10758_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_04018_),
    .Y(_04029_));
 sky130_fd_sc_hd__mux2_1 _10759_ (.A0(_04028_),
    .A1(_04029_),
    .S(_03669_),
    .X(_04030_));
 sky130_fd_sc_hd__and2_1 _10760_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__o21ai_1 _10761_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_04030_),
    .B1(_03997_),
    .Y(_04032_));
 sky130_fd_sc_hd__o221a_1 _10762_ (.A1(_04023_),
    .A2(net463),
    .B1(_04031_),
    .B2(_04032_),
    .C1(_03814_),
    .X(_00493_));
 sky130_fd_sc_hd__inv_2 _10763_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_04033_));
 sky130_fd_sc_hd__buf_2 _10764_ (.A(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__clkbuf_4 _10765_ (.A(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__o21ai_1 _10766_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_04028_),
    .B1(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__a31o_1 _10767_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(_04018_),
    .B1(_04035_),
    .X(_04037_));
 sky130_fd_sc_hd__inv_2 _10768_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .Y(_04038_));
 sky130_fd_sc_hd__a21oi_1 _10769_ (.A1(_04036_),
    .A2(_04037_),
    .B1(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__a31o_1 _10770_ (.A1(_04038_),
    .A2(_04036_),
    .A3(_04037_),
    .B1(_03994_),
    .X(_04040_));
 sky130_fd_sc_hd__o221a_1 _10771_ (.A1(_04023_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_04039_),
    .B2(_04040_),
    .C1(_03814_),
    .X(_00494_));
 sky130_fd_sc_hd__and4_1 _10772_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .D(_04018_),
    .X(_04041_));
 sky130_fd_sc_hd__or3_1 _10773_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C(_04028_),
    .X(_04042_));
 sky130_fd_sc_hd__inv_2 _10774_ (.A(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(_04041_),
    .A1(_04043_),
    .S(_04035_),
    .X(_04044_));
 sky130_fd_sc_hd__xnor2_1 _10776_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_1 _10777_ (.A(_04012_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__o211a_1 _10778_ (.A1(_04011_),
    .A2(net538),
    .B1(_04003_),
    .C1(_04046_),
    .X(_00495_));
 sky130_fd_sc_hd__clkbuf_4 _10779_ (.A(_03993_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_4 _10780_ (.A(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _10781_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_04042_),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_1 _10782_ (.A(_03669_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__a31o_1 _10783_ (.A1(_03669_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_04041_),
    .B1(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__xor2_1 _10784_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(_03999_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(_04053_));
 sky130_fd_sc_hd__o211a_1 _10786_ (.A1(_04048_),
    .A2(_04052_),
    .B1(_04053_),
    .C1(_03780_),
    .X(_00496_));
 sky130_fd_sc_hd__o21a_1 _10787_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_04049_),
    .B1(_04035_),
    .X(_04054_));
 sky130_fd_sc_hd__a31o_1 _10788_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_04041_),
    .B1(_04035_),
    .X(_04055_));
 sky130_fd_sc_hd__or2b_1 _10789_ (.A(_04054_),
    .B_N(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__nor2_1 _10790_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__a21o_1 _10791_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_04056_),
    .B1(_03994_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_4 _10792_ (.A(_02308_),
    .X(_04059_));
 sky130_fd_sc_hd__o221a_1 _10793_ (.A1(_04023_),
    .A2(net422),
    .B1(_04057_),
    .B2(_04058_),
    .C1(_04059_),
    .X(_00497_));
 sky130_fd_sc_hd__a21oi_1 _10794_ (.A1(net651),
    .A2(_04055_),
    .B1(_04054_),
    .Y(_04060_));
 sky130_fd_sc_hd__clkbuf_4 _10795_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_04061_));
 sky130_fd_sc_hd__or2_1 _10796_ (.A(_03999_),
    .B(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_4 _10797_ (.A(_01474_),
    .X(_04063_));
 sky130_fd_sc_hd__o211a_1 _10798_ (.A1(_04048_),
    .A2(_04060_),
    .B1(_04062_),
    .C1(_04063_),
    .X(_00498_));
 sky130_fd_sc_hd__inv_2 _10799_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_04064_));
 sky130_fd_sc_hd__nor2_1 _10800_ (.A(_04064_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_04065_));
 sky130_fd_sc_hd__a21o_1 _10801_ (.A1(_04064_),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_03994_),
    .X(_04066_));
 sky130_fd_sc_hd__o221a_1 _10802_ (.A1(_04023_),
    .A2(net400),
    .B1(_04065_),
    .B2(_04066_),
    .C1(_04059_),
    .X(_00499_));
 sky130_fd_sc_hd__and2b_1 _10803_ (.A_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .X(_04067_));
 sky130_fd_sc_hd__xnor2_1 _10804_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__xnor2_1 _10805_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__xor2_1 _10806_ (.A(_04065_),
    .B(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__or2_1 _10807_ (.A(_04010_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_04071_));
 sky130_fd_sc_hd__o211a_1 _10808_ (.A1(_04048_),
    .A2(_04070_),
    .B1(_04071_),
    .C1(_04063_),
    .X(_00500_));
 sky130_fd_sc_hd__and2_1 _10809_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_04068_),
    .X(_04072_));
 sky130_fd_sc_hd__nor2_1 _10810_ (.A(_04065_),
    .B(_04069_),
    .Y(_04073_));
 sky130_fd_sc_hd__o21ba_1 _10811_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_04074_));
 sky130_fd_sc_hd__xnor2_1 _10812_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__or2_1 _10813_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_04075_),
    .Y(_04077_));
 sky130_fd_sc_hd__and2_1 _10815_ (.A(_04076_),
    .B(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__o21ai_1 _10816_ (.A1(_04072_),
    .A2(_04073_),
    .B1(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__o31a_1 _10817_ (.A1(_04072_),
    .A2(_04073_),
    .A3(_04078_),
    .B1(_03996_),
    .X(_04080_));
 sky130_fd_sc_hd__a22oi_1 _10818_ (.A1(_04047_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_04079_),
    .B2(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__and2b_1 _10819_ (.A_N(_04081_),
    .B(_03118_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _10820_ (.A(_04082_),
    .X(_00501_));
 sky130_fd_sc_hd__o31a_1 _10821_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A3(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1(_04033_),
    .X(_04083_));
 sky130_fd_sc_hd__xnor2_1 _10822_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _10823_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__or2_1 _10824_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_04084_),
    .X(_04086_));
 sky130_fd_sc_hd__and2_1 _10825_ (.A(_04085_),
    .B(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__nand2_1 _10826_ (.A(_04077_),
    .B(_04079_),
    .Y(_04088_));
 sky130_fd_sc_hd__xor2_1 _10827_ (.A(_04087_),
    .B(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_04089_),
    .S(_03996_),
    .X(_04090_));
 sky130_fd_sc_hd__and2_1 _10829_ (.A(_03976_),
    .B(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_04091_),
    .X(_00502_));
 sky130_fd_sc_hd__a21bo_1 _10831_ (.A1(_04077_),
    .A2(_04079_),
    .B1_N(_04087_),
    .X(_04092_));
 sky130_fd_sc_hd__or4_1 _10832_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .C(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .D(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .X(_04093_));
 sky130_fd_sc_hd__nand2_1 _10833_ (.A(_04034_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__xor2_2 _10834_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__xnor2_1 _10835_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__a21oi_1 _10836_ (.A1(_04085_),
    .A2(_04092_),
    .B1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__and3_1 _10837_ (.A(_04085_),
    .B(_04092_),
    .C(_04096_),
    .X(_04098_));
 sky130_fd_sc_hd__o21ai_1 _10838_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04012_),
    .Y(_04099_));
 sky130_fd_sc_hd__o211a_1 _10839_ (.A1(_04011_),
    .A2(net333),
    .B1(_04003_),
    .C1(_04099_),
    .X(_00503_));
 sky130_fd_sc_hd__o21a_1 _10840_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_04093_),
    .B1(_04033_),
    .X(_04100_));
 sky130_fd_sc_hd__xor2_1 _10841_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__or2b_1 _10842_ (.A(_04101_),
    .B_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_04102_));
 sky130_fd_sc_hd__or2b_1 _10843_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B_N(_04101_),
    .X(_04103_));
 sky130_fd_sc_hd__nand2_1 _10844_ (.A(_04102_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__a21oi_1 _10845_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(_04095_),
    .B1(_04097_),
    .Y(_04105_));
 sky130_fd_sc_hd__xor2_1 _10846_ (.A(_04104_),
    .B(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__or2_1 _10847_ (.A(_04010_),
    .B(net543),
    .X(_04107_));
 sky130_fd_sc_hd__o211a_1 _10848_ (.A1(_04048_),
    .A2(_04106_),
    .B1(_04107_),
    .C1(_04063_),
    .X(_00504_));
 sky130_fd_sc_hd__or3_4 _10849_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .C(_04093_),
    .X(_04108_));
 sky130_fd_sc_hd__and2_1 _10850_ (.A(_04034_),
    .B(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__xnor2_1 _10851_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__nand2_1 _10852_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__or2_1 _10853_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_04110_),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _10854_ (.A(_04111_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__a21bo_1 _10855_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .A2(_04095_),
    .B1_N(_04102_),
    .X(_04114_));
 sky130_fd_sc_hd__o21ai_1 _10856_ (.A1(_04097_),
    .A2(_04114_),
    .B1(_04103_),
    .Y(_04115_));
 sky130_fd_sc_hd__xor2_1 _10857_ (.A(_04113_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__mux2_1 _10858_ (.A0(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A1(_04116_),
    .S(_03996_),
    .X(_04117_));
 sky130_fd_sc_hd__and2_1 _10859_ (.A(_03976_),
    .B(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_04118_),
    .X(_00505_));
 sky130_fd_sc_hd__o21a_1 _10861_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_04108_),
    .B1(_04034_),
    .X(_04119_));
 sky130_fd_sc_hd__xor2_1 _10862_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__or2b_1 _10863_ (.A(_04120_),
    .B_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04121_));
 sky130_fd_sc_hd__or2b_1 _10864_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B_N(_04120_),
    .X(_04122_));
 sky130_fd_sc_hd__nand2_1 _10865_ (.A(_04121_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__o21ai_1 _10866_ (.A1(_04113_),
    .A2(_04115_),
    .B1(_04111_),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_1 _10867_ (.A(_04123_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__or2_1 _10868_ (.A(_04010_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04126_));
 sky130_fd_sc_hd__o211a_1 _10869_ (.A1(_04048_),
    .A2(_04125_),
    .B1(_04126_),
    .C1(_04063_),
    .X(_00506_));
 sky130_fd_sc_hd__and2b_1 _10870_ (.A_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_04120_),
    .X(_04127_));
 sky130_fd_sc_hd__a21o_1 _10871_ (.A1(_04111_),
    .A2(_04121_),
    .B1(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__or4bb_1 _10872_ (.A(_04113_),
    .B(_04123_),
    .C_N(_04114_),
    .D_N(_04103_),
    .X(_04129_));
 sky130_fd_sc_hd__or2_1 _10873_ (.A(_04096_),
    .B(_04104_),
    .X(_04130_));
 sky130_fd_sc_hd__a2111o_1 _10874_ (.A1(_04085_),
    .A2(_04092_),
    .B1(_04113_),
    .C1(_04130_),
    .D1(_04123_),
    .X(_04131_));
 sky130_fd_sc_hd__or2_1 _10875_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_04132_));
 sky130_fd_sc_hd__o21ai_1 _10876_ (.A1(_04108_),
    .A2(_04132_),
    .B1(_04035_),
    .Y(_04133_));
 sky130_fd_sc_hd__xor2_1 _10877_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__nand2_1 _10878_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__or2_1 _10879_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04134_),
    .X(_04136_));
 sky130_fd_sc_hd__nand2_1 _10880_ (.A(_04135_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__nand4_1 _10881_ (.A(_04128_),
    .B(_04129_),
    .C(_04131_),
    .D(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__a31o_1 _10882_ (.A1(_04128_),
    .A2(_04129_),
    .A3(_04131_),
    .B1(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__and2_1 _10883_ (.A(_04138_),
    .B(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__or2_1 _10884_ (.A(_04010_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_04141_));
 sky130_fd_sc_hd__o211a_1 _10885_ (.A1(_04048_),
    .A2(_04140_),
    .B1(_04141_),
    .C1(_04063_),
    .X(_00507_));
 sky130_fd_sc_hd__inv_2 _10886_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .Y(_04142_));
 sky130_fd_sc_hd__o31a_2 _10887_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_04108_),
    .A3(_04132_),
    .B1(_04035_),
    .X(_04143_));
 sky130_fd_sc_hd__xor2_4 _10888_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__xnor2_2 _10889_ (.A(_04142_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_1 _10890_ (.A(_04135_),
    .B(_04139_),
    .Y(_04146_));
 sky130_fd_sc_hd__and2_1 _10891_ (.A(_04145_),
    .B(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__o21ai_1 _10892_ (.A1(_04145_),
    .A2(_04146_),
    .B1(_03997_),
    .Y(_04148_));
 sky130_fd_sc_hd__o221a_1 _10893_ (.A1(_04023_),
    .A2(net118),
    .B1(_04147_),
    .B2(_04148_),
    .C1(_04059_),
    .X(_00508_));
 sky130_fd_sc_hd__or3_1 _10894_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .C(_04132_),
    .X(_04149_));
 sky130_fd_sc_hd__or2_1 _10895_ (.A(_04108_),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__and2_1 _10896_ (.A(_04034_),
    .B(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__xnor2_1 _10897_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__nand2_1 _10898_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__or2_1 _10899_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04152_),
    .X(_04154_));
 sky130_fd_sc_hd__nand2_1 _10900_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__o21a_1 _10901_ (.A1(_04142_),
    .A2(_04144_),
    .B1(_04135_),
    .X(_04156_));
 sky130_fd_sc_hd__a21oi_1 _10902_ (.A1(_04142_),
    .A2(_04144_),
    .B1(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__inv_2 _10903_ (.A(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__o21ai_1 _10904_ (.A1(_04139_),
    .A2(_04145_),
    .B1(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__xnor2_1 _10905_ (.A(_04155_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A1(_04160_),
    .S(_03996_),
    .X(_04161_));
 sky130_fd_sc_hd__and2_1 _10907_ (.A(_03976_),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_04162_),
    .X(_00509_));
 sky130_fd_sc_hd__or2b_1 _10909_ (.A(_04155_),
    .B_N(_04159_),
    .X(_04163_));
 sky130_fd_sc_hd__inv_2 _10910_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_04164_));
 sky130_fd_sc_hd__o211a_1 _10911_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_04150_),
    .B1(_04034_),
    .C1(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__a21oi_2 _10912_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B1(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__or3_1 _10913_ (.A(_04164_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .C(_04150_),
    .X(_04167_));
 sky130_fd_sc_hd__a21o_1 _10914_ (.A1(_04166_),
    .A2(_04167_),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_04168_));
 sky130_fd_sc_hd__nand3_1 _10915_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_04166_),
    .C(_04167_),
    .Y(_04169_));
 sky130_fd_sc_hd__and2_1 _10916_ (.A(_04168_),
    .B(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__a21oi_1 _10917_ (.A1(_04153_),
    .A2(_04163_),
    .B1(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__a31o_1 _10918_ (.A1(_04153_),
    .A2(_04163_),
    .A3(_04170_),
    .B1(_03994_),
    .X(_04172_));
 sky130_fd_sc_hd__o221a_1 _10919_ (.A1(_04023_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_04171_),
    .B2(_04172_),
    .C1(_04059_),
    .X(_00510_));
 sky130_fd_sc_hd__or2b_1 _10920_ (.A(_04155_),
    .B_N(_04170_),
    .X(_04173_));
 sky130_fd_sc_hd__or3_1 _10921_ (.A(_04139_),
    .B(_04145_),
    .C(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__or2_1 _10922_ (.A(_04158_),
    .B(_04173_),
    .X(_04175_));
 sky130_fd_sc_hd__or2b_1 _10923_ (.A(_04153_),
    .B_N(_04168_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_4 _10924_ (.A(_04166_),
    .X(_04177_));
 sky130_fd_sc_hd__xnor2_1 _10925_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__a41o_1 _10926_ (.A1(_04169_),
    .A2(_04174_),
    .A3(_04175_),
    .A4(_04176_),
    .B1(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__and4_1 _10927_ (.A(_04169_),
    .B(_04174_),
    .C(_04175_),
    .D(_04176_),
    .X(_04180_));
 sky130_fd_sc_hd__nand2_1 _10928_ (.A(_04178_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__and2_1 _10929_ (.A(_04179_),
    .B(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(_04010_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_04183_));
 sky130_fd_sc_hd__o211a_1 _10931_ (.A1(_04048_),
    .A2(_04182_),
    .B1(_04183_),
    .C1(_04063_),
    .X(_00511_));
 sky130_fd_sc_hd__xnor2_2 _10932_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_04177_),
    .Y(_04184_));
 sky130_fd_sc_hd__a21bo_1 _10933_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_04177_),
    .B1_N(_04179_),
    .X(_04185_));
 sky130_fd_sc_hd__and2_1 _10934_ (.A(_04184_),
    .B(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__o21ai_1 _10935_ (.A1(_04184_),
    .A2(_04185_),
    .B1(_03997_),
    .Y(_04187_));
 sky130_fd_sc_hd__o221a_1 _10936_ (.A1(_04023_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_04186_),
    .B2(_04187_),
    .C1(_04059_),
    .X(_00512_));
 sky130_fd_sc_hd__inv_2 _10937_ (.A(_04177_),
    .Y(_04188_));
 sky130_fd_sc_hd__nor2_1 _10938_ (.A(_03801_),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_1 _10939_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04177_),
    .Y(_04190_));
 sky130_fd_sc_hd__or2_1 _10940_ (.A(_04189_),
    .B(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__nor2_1 _10941_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .Y(_04192_));
 sky130_fd_sc_hd__o22a_1 _10942_ (.A1(_04179_),
    .A2(_04184_),
    .B1(_04192_),
    .B2(_04188_),
    .X(_04193_));
 sky130_fd_sc_hd__nor2_1 _10943_ (.A(_04191_),
    .B(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__and2_1 _10944_ (.A(_04191_),
    .B(_04193_),
    .X(_04195_));
 sky130_fd_sc_hd__nor2_1 _10945_ (.A(_04194_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__or2_1 _10946_ (.A(_04010_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .X(_04197_));
 sky130_fd_sc_hd__o211a_1 _10947_ (.A1(_04048_),
    .A2(_04196_),
    .B1(_04197_),
    .C1(_04063_),
    .X(_00513_));
 sky130_fd_sc_hd__xnor2_1 _10948_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_04177_),
    .Y(_04198_));
 sky130_fd_sc_hd__o21ai_1 _10949_ (.A1(_04189_),
    .A2(_04194_),
    .B1(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__o31a_1 _10950_ (.A1(_04189_),
    .A2(_04194_),
    .A3(_04198_),
    .B1(_03997_),
    .X(_04200_));
 sky130_fd_sc_hd__o21ai_1 _10951_ (.A1(_03997_),
    .A2(net554),
    .B1(_01794_),
    .Y(_04201_));
 sky130_fd_sc_hd__a21oi_1 _10952_ (.A1(_04199_),
    .A2(_04200_),
    .B1(_04201_),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2_1 _10953_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04177_),
    .Y(_04202_));
 sky130_fd_sc_hd__and2_1 _10954_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04177_),
    .X(_04203_));
 sky130_fd_sc_hd__or2_1 _10955_ (.A(_04202_),
    .B(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__or4_1 _10956_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .C(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .D(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_04205_));
 sky130_fd_sc_hd__or3_1 _10957_ (.A(_04184_),
    .B(_04191_),
    .C(_04198_),
    .X(_04206_));
 sky130_fd_sc_hd__o2bb2a_1 _10958_ (.A1_N(_04177_),
    .A2_N(_04205_),
    .B1(_04206_),
    .B2(_04179_),
    .X(_04207_));
 sky130_fd_sc_hd__a21o_1 _10959_ (.A1(_04204_),
    .A2(_04207_),
    .B1(_03993_),
    .X(_04208_));
 sky130_fd_sc_hd__nor2_1 _10960_ (.A(_04204_),
    .B(_04207_),
    .Y(_04209_));
 sky130_fd_sc_hd__a2bb2o_1 _10961_ (.A1_N(_04208_),
    .A2_N(_04209_),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B2(_03993_),
    .X(_04210_));
 sky130_fd_sc_hd__and2_1 _10962_ (.A(_03976_),
    .B(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(_04211_),
    .X(_00515_));
 sky130_fd_sc_hd__xnor2_1 _10964_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_04177_),
    .Y(_04212_));
 sky130_fd_sc_hd__o21ai_1 _10965_ (.A1(_04203_),
    .A2(_04209_),
    .B1(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__o31a_1 _10966_ (.A1(_04203_),
    .A2(_04209_),
    .A3(_04212_),
    .B1(_03997_),
    .X(_04214_));
 sky130_fd_sc_hd__o21ai_1 _10967_ (.A1(_03997_),
    .A2(net642),
    .B1(_01794_),
    .Y(_04215_));
 sky130_fd_sc_hd__a21oi_1 _10968_ (.A1(_04213_),
    .A2(_04214_),
    .B1(_04215_),
    .Y(_00516_));
 sky130_fd_sc_hd__and2_1 _10969_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .X(_04216_));
 sky130_fd_sc_hd__nor2_1 _10970_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .Y(_04217_));
 sky130_fd_sc_hd__o21ai_1 _10971_ (.A1(_04216_),
    .A2(_04217_),
    .B1(_04012_),
    .Y(_04218_));
 sky130_fd_sc_hd__o211a_1 _10972_ (.A1(_04011_),
    .A2(net282),
    .B1(_04003_),
    .C1(_04218_),
    .X(_00517_));
 sky130_fd_sc_hd__buf_4 _10973_ (.A(_03619_),
    .X(_04219_));
 sky130_fd_sc_hd__and2b_1 _10974_ (.A_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .X(_04220_));
 sky130_fd_sc_hd__xnor2_1 _10975_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__xnor2_1 _10976_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__nor2_1 _10977_ (.A(_04216_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__and2_1 _10978_ (.A(_04216_),
    .B(_04222_),
    .X(_04224_));
 sky130_fd_sc_hd__o21ai_1 _10979_ (.A1(_04223_),
    .A2(_04224_),
    .B1(_04012_),
    .Y(_04225_));
 sky130_fd_sc_hd__o211a_1 _10980_ (.A1(_04011_),
    .A2(net419),
    .B1(_04219_),
    .C1(_04225_),
    .X(_00518_));
 sky130_fd_sc_hd__and2b_1 _10981_ (.A_N(_04221_),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_04226_));
 sky130_fd_sc_hd__inv_2 _10982_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_04227_));
 sky130_fd_sc_hd__o21a_1 _10983_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_04034_),
    .X(_04228_));
 sky130_fd_sc_hd__xnor2_1 _10984_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__xnor2_1 _10985_ (.A(_04227_),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__o21bai_2 _10986_ (.A1(_04226_),
    .A2(_04224_),
    .B1_N(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__or3b_1 _10987_ (.A(_04226_),
    .B(_04224_),
    .C_N(_04230_),
    .X(_04232_));
 sky130_fd_sc_hd__inv_2 _10988_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_04233_));
 sky130_fd_sc_hd__nor2_1 _10989_ (.A(_03996_),
    .B(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__a31o_1 _10990_ (.A1(_03996_),
    .A2(_04231_),
    .A3(_04232_),
    .B1(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__and2_1 _10991_ (.A(_03976_),
    .B(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(_04236_),
    .X(_00519_));
 sky130_fd_sc_hd__inv_2 _10993_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_04237_));
 sky130_fd_sc_hd__or2_1 _10994_ (.A(_04227_),
    .B(_04229_),
    .X(_04238_));
 sky130_fd_sc_hd__inv_2 _10995_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_04239_));
 sky130_fd_sc_hd__o31a_1 _10996_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A3(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_04034_),
    .X(_04240_));
 sky130_fd_sc_hd__xnor2_1 _10997_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_1 _10998_ (.A(_04239_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__and2_1 _10999_ (.A(_04239_),
    .B(_04241_),
    .X(_04243_));
 sky130_fd_sc_hd__or2_1 _11000_ (.A(_04242_),
    .B(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__and3_1 _11001_ (.A(_04238_),
    .B(_04231_),
    .C(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__a21oi_1 _11002_ (.A1(_04238_),
    .A2(_04231_),
    .B1(_04244_),
    .Y(_04246_));
 sky130_fd_sc_hd__or3_1 _11003_ (.A(_03993_),
    .B(_04245_),
    .C(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__o21a_1 _11004_ (.A1(_03996_),
    .A2(_04237_),
    .B1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__and2b_1 _11005_ (.A_N(_04248_),
    .B(_03118_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_04249_),
    .X(_00520_));
 sky130_fd_sc_hd__inv_2 _11007_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_04250_));
 sky130_fd_sc_hd__or4_2 _11008_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .C(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .D(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .X(_04251_));
 sky130_fd_sc_hd__nand2_1 _11009_ (.A(_04034_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__xor2_1 _11010_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__or2_1 _11011_ (.A(_04250_),
    .B(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__nand2_1 _11012_ (.A(_04250_),
    .B(_04253_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_1 _11013_ (.A(_04254_),
    .B(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__inv_2 _11014_ (.A(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__o21a_1 _11015_ (.A1(_04242_),
    .A2(_04246_),
    .B1(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__inv_2 _11016_ (.A(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__or3_1 _11017_ (.A(_04242_),
    .B(_04246_),
    .C(_04257_),
    .X(_04260_));
 sky130_fd_sc_hd__a21o_1 _11018_ (.A1(_04259_),
    .A2(_04260_),
    .B1(_04048_),
    .X(_04261_));
 sky130_fd_sc_hd__o211a_1 _11019_ (.A1(_04011_),
    .A2(net571),
    .B1(_04219_),
    .C1(_04261_),
    .X(_00521_));
 sky130_fd_sc_hd__o21a_1 _11020_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_04251_),
    .B1(_04035_),
    .X(_04262_));
 sky130_fd_sc_hd__xor2_1 _11021_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__and2_1 _11022_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__nor2_1 _11023_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_04263_),
    .Y(_04265_));
 sky130_fd_sc_hd__nor2_1 _11024_ (.A(_04264_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__a21oi_1 _11025_ (.A1(_04254_),
    .A2(_04259_),
    .B1(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a31o_1 _11026_ (.A1(_04254_),
    .A2(_04259_),
    .A3(_04266_),
    .B1(_03994_),
    .X(_04268_));
 sky130_fd_sc_hd__o221a_1 _11027_ (.A1(_04023_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B1(_04267_),
    .B2(_04268_),
    .C1(_04059_),
    .X(_00522_));
 sky130_fd_sc_hd__nor3_1 _11028_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .C(_04251_),
    .Y(_04269_));
 sky130_fd_sc_hd__nor2_1 _11029_ (.A(_03669_),
    .B(net115),
    .Y(_04270_));
 sky130_fd_sc_hd__xnor2_2 _11030_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__xnor2_1 _11031_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__a21bo_1 _11032_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(_04263_),
    .B1_N(_04254_),
    .X(_04273_));
 sky130_fd_sc_hd__o21bai_2 _11033_ (.A1(_04258_),
    .A2(_04273_),
    .B1_N(_04265_),
    .Y(_04274_));
 sky130_fd_sc_hd__xnor2_1 _11034_ (.A(_04272_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_04275_),
    .S(_03996_),
    .X(_04276_));
 sky130_fd_sc_hd__and2_1 _11036_ (.A(_03976_),
    .B(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _11037_ (.A(_04277_),
    .X(_00523_));
 sky130_fd_sc_hd__or2_1 _11038_ (.A(_04064_),
    .B(_04271_),
    .X(_04278_));
 sky130_fd_sc_hd__inv_2 _11039_ (.A(_04272_),
    .Y(_04279_));
 sky130_fd_sc_hd__or2_1 _11040_ (.A(_04279_),
    .B(_04274_),
    .X(_04280_));
 sky130_fd_sc_hd__or3_1 _11041_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .C(_04251_),
    .X(_04281_));
 sky130_fd_sc_hd__o21a_1 _11042_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_04281_),
    .B1(_04035_),
    .X(_04282_));
 sky130_fd_sc_hd__xor2_1 _11043_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__nor2_1 _11044_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_1 _11045_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_04283_),
    .Y(_04285_));
 sky130_fd_sc_hd__or2b_1 _11046_ (.A(_04284_),
    .B_N(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__inv_2 _11047_ (.A(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__a21oi_1 _11048_ (.A1(_04278_),
    .A2(_04280_),
    .B1(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__a31o_1 _11049_ (.A1(_04278_),
    .A2(_04280_),
    .A3(_04287_),
    .B1(_04047_),
    .X(_04289_));
 sky130_fd_sc_hd__o221a_1 _11050_ (.A1(_04023_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B1(_04288_),
    .B2(_04289_),
    .C1(_04059_),
    .X(_00524_));
 sky130_fd_sc_hd__o21a_1 _11051_ (.A1(_04278_),
    .A2(_04284_),
    .B1(_04285_),
    .X(_04290_));
 sky130_fd_sc_hd__o21a_1 _11052_ (.A1(_04280_),
    .A2(_04286_),
    .B1(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__inv_2 _11053_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_04292_));
 sky130_fd_sc_hd__a21oi_1 _11054_ (.A1(_04192_),
    .A2(net115),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_04293_));
 sky130_fd_sc_hd__xnor2_1 _11055_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__or2_1 _11056_ (.A(_04292_),
    .B(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__nand2_1 _11057_ (.A(_04292_),
    .B(_04294_),
    .Y(_04296_));
 sky130_fd_sc_hd__nand2_1 _11058_ (.A(_04295_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2_1 _11059_ (.A(_04291_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__or2_1 _11060_ (.A(_04291_),
    .B(_04297_),
    .X(_04299_));
 sky130_fd_sc_hd__a21o_1 _11061_ (.A1(_04298_),
    .A2(_04299_),
    .B1(_03994_),
    .X(_04300_));
 sky130_fd_sc_hd__o211a_1 _11062_ (.A1(_04011_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_04219_),
    .C1(_04300_),
    .X(_00525_));
 sky130_fd_sc_hd__a31o_1 _11063_ (.A1(_03801_),
    .A2(_04192_),
    .A3(net115),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_04301_));
 sky130_fd_sc_hd__xnor2_1 _11064_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _11065_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__or2_1 _11066_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__nand2_1 _11067_ (.A(_04303_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__o21ai_1 _11068_ (.A1(_04291_),
    .A2(_04297_),
    .B1(_04295_),
    .Y(_04306_));
 sky130_fd_sc_hd__nor2_1 _11069_ (.A(_04305_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21o_1 _11070_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_03994_),
    .X(_04308_));
 sky130_fd_sc_hd__o221a_1 _11071_ (.A1(_04012_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_04307_),
    .B2(_04308_),
    .C1(_04059_),
    .X(_00526_));
 sky130_fd_sc_hd__a21bo_1 _11072_ (.A1(_04295_),
    .A2(_04303_),
    .B1_N(_04304_),
    .X(_04309_));
 sky130_fd_sc_hd__o31ai_2 _11073_ (.A1(_04279_),
    .A2(_04274_),
    .A3(_04286_),
    .B1(_04290_),
    .Y(_04310_));
 sky130_fd_sc_hd__nor2_1 _11074_ (.A(_04297_),
    .B(_04305_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _11075_ (.A(_04310_),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__or2_1 _11076_ (.A(_04205_),
    .B(_04281_),
    .X(_04313_));
 sky130_fd_sc_hd__nand2_1 _11077_ (.A(_04035_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__xor2_1 _11078_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__inv_2 _11079_ (.A(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _11080_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__or2_1 _11081_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04316_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _11082_ (.A(_04317_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a21o_1 _11083_ (.A1(_04309_),
    .A2(_04312_),
    .B1(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__a31oi_1 _11084_ (.A1(_04319_),
    .A2(_04309_),
    .A3(_04312_),
    .B1(_03993_),
    .Y(_04321_));
 sky130_fd_sc_hd__a22o_1 _11085_ (.A1(_04047_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_04320_),
    .B2(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__and2_1 _11086_ (.A(_03976_),
    .B(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _11087_ (.A(_04323_),
    .X(_00527_));
 sky130_fd_sc_hd__o21a_1 _11088_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(_04313_),
    .B1(_04034_),
    .X(_04324_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(_04324_),
    .A1(_03669_),
    .S(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_04325_));
 sky130_fd_sc_hd__and4bb_1 _11090_ (.A_N(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B_N(_04205_),
    .C(net115),
    .D(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_04326_));
 sky130_fd_sc_hd__or3_1 _11091_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04325_),
    .C(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__o21ai_2 _11092_ (.A1(_04325_),
    .A2(_04326_),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .Y(_04328_));
 sky130_fd_sc_hd__and2_1 _11093_ (.A(_04327_),
    .B(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__a21oi_1 _11094_ (.A1(_04317_),
    .A2(_04320_),
    .B1(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__a31o_1 _11095_ (.A1(_04317_),
    .A2(_04320_),
    .A3(_04329_),
    .B1(_04047_),
    .X(_04331_));
 sky130_fd_sc_hd__o221a_1 _11096_ (.A1(_04012_),
    .A2(net621),
    .B1(_04330_),
    .B2(_04331_),
    .C1(_04059_),
    .X(_00528_));
 sky130_fd_sc_hd__and3b_1 _11097_ (.A_N(_04319_),
    .B(_04311_),
    .C(_04329_),
    .X(_04332_));
 sky130_fd_sc_hd__and4bb_1 _11098_ (.A_N(_04319_),
    .B_N(_04309_),
    .C(_04327_),
    .D(_04328_),
    .X(_04333_));
 sky130_fd_sc_hd__inv_2 _11099_ (.A(_04328_),
    .Y(_04334_));
 sky130_fd_sc_hd__a31o_1 _11100_ (.A1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_04316_),
    .A3(_04327_),
    .B1(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__a211o_1 _11101_ (.A1(_04310_),
    .A2(_04332_),
    .B1(_04333_),
    .C1(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__or2_1 _11102_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_04325_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_4 _11103_ (.A(_04325_),
    .X(_04338_));
 sky130_fd_sc_hd__nand2_1 _11104_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__and2_1 _11105_ (.A(_04337_),
    .B(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__nand2_1 _11106_ (.A(_04336_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__or2_1 _11107_ (.A(_04336_),
    .B(_04340_),
    .X(_04342_));
 sky130_fd_sc_hd__and2_1 _11108_ (.A(_04341_),
    .B(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__or2_1 _11109_ (.A(_04010_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_04344_));
 sky130_fd_sc_hd__o211a_1 _11110_ (.A1(_04048_),
    .A2(_04343_),
    .B1(_04344_),
    .C1(_04063_),
    .X(_00529_));
 sky130_fd_sc_hd__xor2_1 _11111_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_04338_),
    .X(_04345_));
 sky130_fd_sc_hd__a21oi_1 _11112_ (.A1(_04339_),
    .A2(_04341_),
    .B1(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__a31o_1 _11113_ (.A1(_04339_),
    .A2(_04341_),
    .A3(_04345_),
    .B1(_04047_),
    .X(_04347_));
 sky130_fd_sc_hd__o221a_1 _11114_ (.A1(_04012_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_04346_),
    .B2(_04347_),
    .C1(_04059_),
    .X(_00530_));
 sky130_fd_sc_hd__or2_1 _11115_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_04338_),
    .X(_04348_));
 sky130_fd_sc_hd__nand2_1 _11116_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_04338_),
    .Y(_04349_));
 sky130_fd_sc_hd__and2_1 _11117_ (.A(_04348_),
    .B(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__and2_1 _11118_ (.A(_04340_),
    .B(_04345_),
    .X(_04351_));
 sky130_fd_sc_hd__a22o_1 _11119_ (.A1(_04132_),
    .A2(_04338_),
    .B1(_04336_),
    .B2(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__nand2_1 _11120_ (.A(_04350_),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__o21a_1 _11121_ (.A1(_04350_),
    .A2(_04352_),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04354_));
 sky130_fd_sc_hd__a22o_1 _11122_ (.A1(_04047_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_04353_),
    .B2(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__and2_1 _11123_ (.A(_03976_),
    .B(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _11124_ (.A(_04356_),
    .X(_00531_));
 sky130_fd_sc_hd__xor2_2 _11125_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_04338_),
    .X(_04357_));
 sky130_fd_sc_hd__a21oi_1 _11126_ (.A1(_04349_),
    .A2(_04353_),
    .B1(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__a31o_1 _11127_ (.A1(_04349_),
    .A2(_04353_),
    .A3(_04357_),
    .B1(_04047_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_4 _11128_ (.A(_02308_),
    .X(_04360_));
 sky130_fd_sc_hd__o221a_1 _11129_ (.A1(_04012_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_04358_),
    .B2(_04359_),
    .C1(_04360_),
    .X(_00532_));
 sky130_fd_sc_hd__and4_1 _11130_ (.A(_04336_),
    .B(_04350_),
    .C(_04351_),
    .D(_04357_),
    .X(_04361_));
 sky130_fd_sc_hd__and2_1 _11131_ (.A(_04149_),
    .B(_04338_),
    .X(_04362_));
 sky130_fd_sc_hd__or2_1 _11132_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04338_),
    .X(_04363_));
 sky130_fd_sc_hd__nand2_1 _11133_ (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04338_),
    .Y(_04364_));
 sky130_fd_sc_hd__and2_1 _11134_ (.A(_04363_),
    .B(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__o21ai_2 _11135_ (.A1(_04361_),
    .A2(_04362_),
    .B1(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__o31a_1 _11136_ (.A1(_04365_),
    .A2(_04361_),
    .A3(_04362_),
    .B1(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04367_));
 sky130_fd_sc_hd__a22o_1 _11137_ (.A1(_04047_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B1(_04366_),
    .B2(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__and2_1 _11138_ (.A(_03976_),
    .B(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _11139_ (.A(_04369_),
    .X(_00533_));
 sky130_fd_sc_hd__xnor2_1 _11140_ (.A(_04164_),
    .B(_04338_),
    .Y(_04370_));
 sky130_fd_sc_hd__a21oi_1 _11141_ (.A1(_04364_),
    .A2(_04366_),
    .B1(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__a31o_1 _11142_ (.A1(_04364_),
    .A2(_04366_),
    .A3(_04370_),
    .B1(_04047_),
    .X(_04372_));
 sky130_fd_sc_hd__o221a_1 _11143_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_04011_),
    .B1(_04371_),
    .B2(_04372_),
    .C1(_04360_),
    .X(_00534_));
 sky130_fd_sc_hd__and2_1 _11144_ (.A(_03997_),
    .B(_02310_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _11145_ (.A(_04373_),
    .X(_00535_));
 sky130_fd_sc_hd__inv_2 _11146_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_04374_));
 sky130_fd_sc_hd__clkbuf_4 _11147_ (.A(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_4 _11148_ (.A(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_4 _11149_ (.A(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_4 _11150_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_2 _11151_ (.A(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__or2_1 _11152_ (.A(net143),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__o211a_1 _11153_ (.A1(_04377_),
    .A2(net157),
    .B1(_04219_),
    .C1(_04380_),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _11154_ (.A(net128),
    .B(_04379_),
    .X(_04381_));
 sky130_fd_sc_hd__o211a_1 _11155_ (.A1(_04377_),
    .A2(net251),
    .B1(_04219_),
    .C1(_04381_),
    .X(_00537_));
 sky130_fd_sc_hd__or2_1 _11156_ (.A(net122),
    .B(_04379_),
    .X(_04382_));
 sky130_fd_sc_hd__o211a_1 _11157_ (.A1(_04377_),
    .A2(net223),
    .B1(_04219_),
    .C1(_04382_),
    .X(_00538_));
 sky130_fd_sc_hd__or2_1 _11158_ (.A(net151),
    .B(_04379_),
    .X(_04383_));
 sky130_fd_sc_hd__o211a_1 _11159_ (.A1(_04377_),
    .A2(net175),
    .B1(_04219_),
    .C1(_04383_),
    .X(_00539_));
 sky130_fd_sc_hd__or2_1 _11160_ (.A(net166),
    .B(_04379_),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _11161_ (.A1(_04377_),
    .A2(net222),
    .B1(_04219_),
    .C1(_04384_),
    .X(_00540_));
 sky130_fd_sc_hd__or2_1 _11162_ (.A(net134),
    .B(_04379_),
    .X(_04385_));
 sky130_fd_sc_hd__o211a_1 _11163_ (.A1(_04377_),
    .A2(net261),
    .B1(_04219_),
    .C1(_04385_),
    .X(_00541_));
 sky130_fd_sc_hd__or2_1 _11164_ (.A(net138),
    .B(_04379_),
    .X(_04386_));
 sky130_fd_sc_hd__o211a_1 _11165_ (.A1(_04377_),
    .A2(net260),
    .B1(_04219_),
    .C1(_04386_),
    .X(_00542_));
 sky130_fd_sc_hd__clkbuf_4 _11166_ (.A(_03619_),
    .X(_04387_));
 sky130_fd_sc_hd__or2_1 _11167_ (.A(net161),
    .B(_04379_),
    .X(_04388_));
 sky130_fd_sc_hd__o211a_1 _11168_ (.A1(_04377_),
    .A2(net276),
    .B1(_04387_),
    .C1(_04388_),
    .X(_00543_));
 sky130_fd_sc_hd__or2_1 _11169_ (.A(_04379_),
    .B(net274),
    .X(_04389_));
 sky130_fd_sc_hd__o211a_1 _11170_ (.A1(_04377_),
    .A2(net290),
    .B1(_04387_),
    .C1(_04389_),
    .X(_00544_));
 sky130_fd_sc_hd__clkbuf_4 _11171_ (.A(_04378_),
    .X(_04390_));
 sky130_fd_sc_hd__buf_4 _11172_ (.A(_04378_),
    .X(_04391_));
 sky130_fd_sc_hd__nand2_1 _11173_ (.A(_04391_),
    .B(net285),
    .Y(_04392_));
 sky130_fd_sc_hd__o211a_1 _11174_ (.A1(_04390_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B1(_04387_),
    .C1(_04392_),
    .X(_00545_));
 sky130_fd_sc_hd__nand2_1 _11175_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_04393_));
 sky130_fd_sc_hd__or2_1 _11176_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(_04394_));
 sky130_fd_sc_hd__a21oi_2 _11177_ (.A1(_04393_),
    .A2(_04394_),
    .B1(_04061_),
    .Y(_04395_));
 sky130_fd_sc_hd__buf_4 _11178_ (.A(_04375_),
    .X(_04396_));
 sky130_fd_sc_hd__a31o_1 _11179_ (.A1(_04061_),
    .A2(_04393_),
    .A3(_04394_),
    .B1(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__o221a_1 _11180_ (.A1(_04390_),
    .A2(net506),
    .B1(_04395_),
    .B2(_04397_),
    .C1(_04360_),
    .X(_00546_));
 sky130_fd_sc_hd__and3_1 _11181_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(_04398_));
 sky130_fd_sc_hd__a21oi_1 _11182_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_04399_));
 sky130_fd_sc_hd__or2_1 _11183_ (.A(_04398_),
    .B(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__nor2_1 _11184_ (.A(_04395_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__a21o_1 _11185_ (.A1(_04395_),
    .A2(_04400_),
    .B1(_04376_),
    .X(_04402_));
 sky130_fd_sc_hd__o221a_1 _11186_ (.A1(_04390_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_04401_),
    .B2(_04402_),
    .C1(_04360_),
    .X(_00547_));
 sky130_fd_sc_hd__nand2_1 _11187_ (.A(_04061_),
    .B(_04398_),
    .Y(_04403_));
 sky130_fd_sc_hd__o31a_1 _11188_ (.A1(_04061_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A3(_04394_),
    .B1(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__and2_1 _11189_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__o21ai_1 _11190_ (.A1(net622),
    .A2(_04404_),
    .B1(_04391_),
    .Y(_04406_));
 sky130_fd_sc_hd__o221a_1 _11191_ (.A1(_04390_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_04405_),
    .B2(_04406_),
    .C1(_04360_),
    .X(_00548_));
 sky130_fd_sc_hd__or3_1 _11192_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(_04394_),
    .X(_04407_));
 sky130_fd_sc_hd__nand2_1 _11193_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_04398_),
    .Y(_04408_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(_04407_),
    .A1(_04408_),
    .S(_04061_),
    .X(_04409_));
 sky130_fd_sc_hd__and2_1 _11195_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__o21ai_1 _11196_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_04409_),
    .B1(_04391_),
    .Y(_04411_));
 sky130_fd_sc_hd__o221a_1 _11197_ (.A1(_04390_),
    .A2(net460),
    .B1(_04410_),
    .B2(_04411_),
    .C1(_04360_),
    .X(_00549_));
 sky130_fd_sc_hd__inv_2 _11198_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_04412_));
 sky130_fd_sc_hd__buf_2 _11199_ (.A(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_4 _11200_ (.A(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__o21ai_1 _11201_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_04407_),
    .B1(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__a31o_1 _11202_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A3(_04398_),
    .B1(_04414_),
    .X(_04416_));
 sky130_fd_sc_hd__inv_2 _11203_ (.A(net463),
    .Y(_04417_));
 sky130_fd_sc_hd__a21oi_1 _11204_ (.A1(_04415_),
    .A2(_04416_),
    .B1(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__a31o_1 _11205_ (.A1(_04417_),
    .A2(_04415_),
    .A3(_04416_),
    .B1(_04396_),
    .X(_04419_));
 sky130_fd_sc_hd__o221a_1 _11206_ (.A1(_04390_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_04418_),
    .B2(_04419_),
    .C1(_04360_),
    .X(_00550_));
 sky130_fd_sc_hd__and4_1 _11207_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .D(_04398_),
    .X(_04420_));
 sky130_fd_sc_hd__or3_1 _11208_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_04407_),
    .X(_04421_));
 sky130_fd_sc_hd__inv_2 _11209_ (.A(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(_04420_),
    .A1(_04422_),
    .S(_04414_),
    .X(_04423_));
 sky130_fd_sc_hd__xnor2_1 _11211_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__nand2_1 _11212_ (.A(_04391_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__o211a_1 _11213_ (.A1(_04390_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_04387_),
    .C1(_04425_),
    .X(_00551_));
 sky130_fd_sc_hd__nand2_1 _11214_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_04420_),
    .Y(_04426_));
 sky130_fd_sc_hd__or2_1 _11215_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_04421_),
    .X(_04427_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(_04426_),
    .A1(_04427_),
    .S(_04414_),
    .X(_04428_));
 sky130_fd_sc_hd__o21ai_1 _11217_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_04428_),
    .B1(_04378_),
    .Y(_04429_));
 sky130_fd_sc_hd__a21o_1 _11218_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_04428_),
    .B1(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__o211a_1 _11219_ (.A1(_04390_),
    .A2(net359),
    .B1(_04387_),
    .C1(_04430_),
    .X(_00552_));
 sky130_fd_sc_hd__buf_4 _11220_ (.A(_04378_),
    .X(_04431_));
 sky130_fd_sc_hd__or2_1 _11221_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_04427_),
    .X(_04432_));
 sky130_fd_sc_hd__a31o_1 _11222_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A3(_04420_),
    .B1(_04414_),
    .X(_04433_));
 sky130_fd_sc_hd__a21bo_1 _11223_ (.A1(_04414_),
    .A2(_04432_),
    .B1_N(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__nor2_1 _11224_ (.A(net387),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a21o_1 _11225_ (.A1(net387),
    .A2(_04434_),
    .B1(_04376_),
    .X(_04436_));
 sky130_fd_sc_hd__o221a_1 _11226_ (.A1(_04431_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_04435_),
    .B2(_04436_),
    .C1(_04360_),
    .X(_00553_));
 sky130_fd_sc_hd__o21a_1 _11227_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_04432_),
    .B1(_04414_),
    .X(_04437_));
 sky130_fd_sc_hd__a41o_1 _11228_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A4(_04420_),
    .B1(_04414_),
    .X(_04438_));
 sky130_fd_sc_hd__or2b_1 _11229_ (.A(_04437_),
    .B_N(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__xnor2_1 _11230_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__or2_1 _11231_ (.A(_04379_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_04441_));
 sky130_fd_sc_hd__o211a_1 _11232_ (.A1(_04377_),
    .A2(_04440_),
    .B1(_04441_),
    .C1(_04063_),
    .X(_00554_));
 sky130_fd_sc_hd__clkbuf_4 _11233_ (.A(_04376_),
    .X(_04442_));
 sky130_fd_sc_hd__a21oi_1 _11234_ (.A1(net422),
    .A2(_04438_),
    .B1(_04437_),
    .Y(_04443_));
 sky130_fd_sc_hd__clkbuf_2 _11235_ (.A(_04378_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_4 _11236_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_04445_));
 sky130_fd_sc_hd__or2_1 _11237_ (.A(_04444_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__o211a_1 _11238_ (.A1(_04442_),
    .A2(_04443_),
    .B1(_04446_),
    .C1(_04063_),
    .X(_00555_));
 sky130_fd_sc_hd__inv_2 _11239_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .Y(_04447_));
 sky130_fd_sc_hd__nor2_1 _11240_ (.A(_04447_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_04448_));
 sky130_fd_sc_hd__a21o_1 _11241_ (.A1(_04447_),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_04376_),
    .X(_04449_));
 sky130_fd_sc_hd__o221a_1 _11242_ (.A1(_04431_),
    .A2(net540),
    .B1(_04448_),
    .B2(_04449_),
    .C1(_04360_),
    .X(_00556_));
 sky130_fd_sc_hd__and2b_1 _11243_ (.A_N(_04061_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_04450_));
 sky130_fd_sc_hd__xnor2_1 _11244_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__xnor2_1 _11245_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__xor2_1 _11246_ (.A(_04448_),
    .B(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__or2_1 _11247_ (.A(_04444_),
    .B(net583),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_8 _11248_ (.A(_01251_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_4 _11249_ (.A(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__o211a_1 _11250_ (.A1(_04442_),
    .A2(_04453_),
    .B1(_04454_),
    .C1(_04456_),
    .X(_00557_));
 sky130_fd_sc_hd__and2_1 _11251_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_04451_),
    .X(_04457_));
 sky130_fd_sc_hd__nor2_1 _11252_ (.A(_04448_),
    .B(_04452_),
    .Y(_04458_));
 sky130_fd_sc_hd__o21ba_1 _11253_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B1_N(_04061_),
    .X(_04459_));
 sky130_fd_sc_hd__xnor2_1 _11254_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__or2_1 _11255_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__nand2_1 _11256_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_04460_),
    .Y(_04462_));
 sky130_fd_sc_hd__and2_1 _11257_ (.A(_04461_),
    .B(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__o21ai_2 _11258_ (.A1(_04457_),
    .A2(_04458_),
    .B1(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__o31a_1 _11259_ (.A1(_04457_),
    .A2(_04458_),
    .A3(_04463_),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04465_));
 sky130_fd_sc_hd__a22oi_1 _11260_ (.A1(_04396_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_04464_),
    .B2(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__and2b_1 _11261_ (.A_N(_04466_),
    .B(_03118_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _11262_ (.A(_04467_),
    .X(_00558_));
 sky130_fd_sc_hd__clkbuf_4 _11263_ (.A(_01252_),
    .X(_04468_));
 sky130_fd_sc_hd__o31a_1 _11264_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A3(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B1(_04412_),
    .X(_04469_));
 sky130_fd_sc_hd__xnor2_1 _11265_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand2_1 _11266_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__or2_1 _11267_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_04470_),
    .X(_04472_));
 sky130_fd_sc_hd__and2_1 _11268_ (.A(_04471_),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__nand2_1 _11269_ (.A(_04462_),
    .B(_04464_),
    .Y(_04474_));
 sky130_fd_sc_hd__xor2_1 _11270_ (.A(_04473_),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__mux2_1 _11271_ (.A0(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_04475_),
    .S(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04476_));
 sky130_fd_sc_hd__and2_1 _11272_ (.A(_04468_),
    .B(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _11273_ (.A(_04477_),
    .X(_00559_));
 sky130_fd_sc_hd__inv_2 _11274_ (.A(_04471_),
    .Y(_04478_));
 sky130_fd_sc_hd__a21boi_2 _11275_ (.A1(_04462_),
    .A2(_04464_),
    .B1_N(_04473_),
    .Y(_04479_));
 sky130_fd_sc_hd__nor2_1 _11276_ (.A(_04478_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__or4_2 _11277_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .C(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .D(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_04481_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(_04413_),
    .B(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__xor2_1 _11279_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__and2_1 _11280_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__nor2_1 _11281_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_04483_),
    .Y(_04485_));
 sky130_fd_sc_hd__or2_1 _11282_ (.A(_04484_),
    .B(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__xor2_1 _11283_ (.A(_04480_),
    .B(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__or2_1 _11284_ (.A(_04444_),
    .B(net491),
    .X(_04488_));
 sky130_fd_sc_hd__o211a_1 _11285_ (.A1(_04442_),
    .A2(_04487_),
    .B1(_04488_),
    .C1(_04456_),
    .X(_00560_));
 sky130_fd_sc_hd__o21a_1 _11286_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(_04481_),
    .B1(_04413_),
    .X(_04489_));
 sky130_fd_sc_hd__xor2_1 _11287_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__and2b_1 _11288_ (.A_N(_04490_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_04491_));
 sky130_fd_sc_hd__or2b_1 _11289_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B_N(_04490_),
    .X(_04492_));
 sky130_fd_sc_hd__or2b_1 _11290_ (.A(_04491_),
    .B_N(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__o21bai_1 _11291_ (.A1(_04480_),
    .A2(_04486_),
    .B1_N(_04484_),
    .Y(_04494_));
 sky130_fd_sc_hd__xnor2_1 _11292_ (.A(_04493_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__or2_1 _11293_ (.A(_04444_),
    .B(net479),
    .X(_04496_));
 sky130_fd_sc_hd__o211a_1 _11294_ (.A1(_04442_),
    .A2(_04495_),
    .B1(_04496_),
    .C1(_04456_),
    .X(_00561_));
 sky130_fd_sc_hd__nor2_1 _11295_ (.A(_04486_),
    .B(_04493_),
    .Y(_04497_));
 sky130_fd_sc_hd__o21a_1 _11296_ (.A1(_04478_),
    .A2(_04479_),
    .B1(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__o21a_1 _11297_ (.A1(_04484_),
    .A2(_04491_),
    .B1(_04492_),
    .X(_04499_));
 sky130_fd_sc_hd__or3_1 _11298_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .C(_04481_),
    .X(_04500_));
 sky130_fd_sc_hd__and2_1 _11299_ (.A(_04413_),
    .B(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__xnor2_1 _11300_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2_1 _11301_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__or2_1 _11302_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_04502_),
    .X(_04504_));
 sky130_fd_sc_hd__and2_1 _11303_ (.A(_04503_),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__o21ai_1 _11304_ (.A1(_04498_),
    .A2(_04499_),
    .B1(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__o31a_1 _11305_ (.A1(_04505_),
    .A2(_04498_),
    .A3(_04499_),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04507_));
 sky130_fd_sc_hd__a22o_1 _11306_ (.A1(_04375_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_04506_),
    .B2(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__and2_1 _11307_ (.A(_04468_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(_04509_),
    .X(_00562_));
 sky130_fd_sc_hd__o21a_1 _11309_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_04500_),
    .B1(_04413_),
    .X(_04510_));
 sky130_fd_sc_hd__xor2_1 _11310_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__and2b_1 _11311_ (.A_N(_04511_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04512_));
 sky130_fd_sc_hd__and2b_1 _11312_ (.A_N(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_04511_),
    .X(_04513_));
 sky130_fd_sc_hd__nor2_1 _11313_ (.A(_04512_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__a21oi_1 _11314_ (.A1(_04503_),
    .A2(_04506_),
    .B1(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__a31o_1 _11315_ (.A1(_04503_),
    .A2(_04506_),
    .A3(_04514_),
    .B1(_04396_),
    .X(_04516_));
 sky130_fd_sc_hd__o221a_1 _11316_ (.A1(_04431_),
    .A2(net544),
    .B1(_04515_),
    .B2(_04516_),
    .C1(_04360_),
    .X(_00563_));
 sky130_fd_sc_hd__or2_1 _11317_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_04517_));
 sky130_fd_sc_hd__or4_4 _11318_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .C(_04481_),
    .D(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__and2_1 _11319_ (.A(_04413_),
    .B(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_1 _11320_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _11321_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__or2_1 _11322_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04520_),
    .X(_04522_));
 sky130_fd_sc_hd__and2_1 _11323_ (.A(_04521_),
    .B(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__or2b_1 _11324_ (.A(_04511_),
    .B_N(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_1 _11325_ (.A1(_04503_),
    .A2(_04524_),
    .B1(_04513_),
    .Y(_04525_));
 sky130_fd_sc_hd__a31o_1 _11326_ (.A1(_04505_),
    .A2(_04499_),
    .A3(_04514_),
    .B1(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__o2111a_1 _11327_ (.A1(_04478_),
    .A2(_04479_),
    .B1(_04505_),
    .C1(_04497_),
    .D1(_04514_),
    .X(_04527_));
 sky130_fd_sc_hd__or3_1 _11328_ (.A(_04523_),
    .B(_04526_),
    .C(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__o21a_1 _11329_ (.A1(_04526_),
    .A2(_04527_),
    .B1(_04523_),
    .X(_04529_));
 sky130_fd_sc_hd__inv_2 _11330_ (.A(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_04528_),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__or2_1 _11332_ (.A(_04444_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_04532_));
 sky130_fd_sc_hd__o211a_1 _11333_ (.A1(_04442_),
    .A2(_04531_),
    .B1(_04532_),
    .C1(_04456_),
    .X(_00564_));
 sky130_fd_sc_hd__o21a_1 _11334_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(_04518_),
    .B1(_04414_),
    .X(_04533_));
 sky130_fd_sc_hd__xor2_2 _11335_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__xnor2_2 _11336_ (.A(net119),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__a21oi_1 _11337_ (.A1(_04521_),
    .A2(_04530_),
    .B1(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__a31o_1 _11338_ (.A1(_04521_),
    .A2(_04530_),
    .A3(_04535_),
    .B1(_04396_),
    .X(_04537_));
 sky130_fd_sc_hd__buf_4 _11339_ (.A(_01251_),
    .X(_04538_));
 sky130_fd_sc_hd__buf_4 _11340_ (.A(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__o221a_1 _11341_ (.A1(_04431_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_04536_),
    .B2(_04537_),
    .C1(_04539_),
    .X(_00565_));
 sky130_fd_sc_hd__inv_2 _11342_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .Y(_04540_));
 sky130_fd_sc_hd__nor3_1 _11343_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .C(_04518_),
    .Y(_04541_));
 sky130_fd_sc_hd__inv_2 _11344_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_04542_));
 sky130_fd_sc_hd__o31a_1 _11345_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A3(_04518_),
    .B1(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__mux2_1 _11346_ (.A0(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A1(_04543_),
    .S(_04413_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_2 _11347_ (.A(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__a21o_1 _11348_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_04541_),
    .B1(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__nor2_1 _11349_ (.A(_04540_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__and2_1 _11350_ (.A(_04540_),
    .B(_04546_),
    .X(_04548_));
 sky130_fd_sc_hd__or2_1 _11351_ (.A(_04547_),
    .B(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__inv_2 _11352_ (.A(net119),
    .Y(_04550_));
 sky130_fd_sc_hd__o2bb2a_1 _11353_ (.A1_N(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2_N(_04520_),
    .B1(_04534_),
    .B2(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__a21oi_1 _11354_ (.A1(_04550_),
    .A2(_04534_),
    .B1(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a21oi_1 _11355_ (.A1(_04529_),
    .A2(_04535_),
    .B1(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__xor2_1 _11356_ (.A(_04549_),
    .B(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__mux2_1 _11357_ (.A0(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A1(_04554_),
    .S(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04555_));
 sky130_fd_sc_hd__and2_1 _11358_ (.A(_04468_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _11359_ (.A(_04556_),
    .X(_00566_));
 sky130_fd_sc_hd__clkbuf_4 _11360_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_04557_));
 sky130_fd_sc_hd__xnor2_1 _11361_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_04545_),
    .Y(_04558_));
 sky130_fd_sc_hd__o21ba_1 _11362_ (.A1(_04549_),
    .A2(_04553_),
    .B1_N(_04547_),
    .X(_04559_));
 sky130_fd_sc_hd__and2_1 _11363_ (.A(_04558_),
    .B(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__o21ai_1 _11364_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04391_),
    .Y(_04561_));
 sky130_fd_sc_hd__o221a_1 _11365_ (.A1(_04431_),
    .A2(_04557_),
    .B1(_04560_),
    .B2(_04561_),
    .C1(_04539_),
    .X(_00567_));
 sky130_fd_sc_hd__and2b_1 _11366_ (.A_N(_04549_),
    .B(_04558_),
    .X(_04562_));
 sky130_fd_sc_hd__and3_1 _11367_ (.A(_04529_),
    .B(_04535_),
    .C(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__or2_1 _11368_ (.A(_04061_),
    .B(_04543_),
    .X(_04564_));
 sky130_fd_sc_hd__o21ai_4 _11369_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_04414_),
    .B1(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__a221o_1 _11370_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_04565_),
    .B1(_04552_),
    .B2(_04562_),
    .C1(_04547_),
    .X(_04566_));
 sky130_fd_sc_hd__or2_1 _11371_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__nand2_1 _11372_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04565_),
    .Y(_04568_));
 sky130_fd_sc_hd__and2_1 _11373_ (.A(_04567_),
    .B(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__o21ai_2 _11374_ (.A1(_04563_),
    .A2(_04566_),
    .B1(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__or3_1 _11375_ (.A(_04569_),
    .B(_04563_),
    .C(_04566_),
    .X(_04571_));
 sky130_fd_sc_hd__and2_1 _11376_ (.A(_04570_),
    .B(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__or2_1 _11377_ (.A(_04444_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_04573_));
 sky130_fd_sc_hd__o211a_1 _11378_ (.A1(_04442_),
    .A2(_04572_),
    .B1(_04573_),
    .C1(_04456_),
    .X(_00568_));
 sky130_fd_sc_hd__xnor2_1 _11379_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_04545_),
    .Y(_04574_));
 sky130_fd_sc_hd__a21oi_1 _11380_ (.A1(_04568_),
    .A2(_04570_),
    .B1(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__a31o_1 _11381_ (.A1(_04568_),
    .A2(_04570_),
    .A3(_04574_),
    .B1(_04396_),
    .X(_04576_));
 sky130_fd_sc_hd__o221a_1 _11382_ (.A1(_04431_),
    .A2(net556),
    .B1(_04575_),
    .B2(_04576_),
    .C1(_04539_),
    .X(_00569_));
 sky130_fd_sc_hd__o21ba_1 _11383_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_04565_),
    .B1_N(_04570_),
    .X(_04577_));
 sky130_fd_sc_hd__o21a_1 _11384_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_04565_),
    .X(_04578_));
 sky130_fd_sc_hd__nand2_1 _11385_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04565_),
    .Y(_04579_));
 sky130_fd_sc_hd__or2_1 _11386_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04565_),
    .X(_04580_));
 sky130_fd_sc_hd__and2_1 _11387_ (.A(_04579_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__o21ai_1 _11388_ (.A1(_04577_),
    .A2(_04578_),
    .B1(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__o31a_1 _11389_ (.A1(_04581_),
    .A2(_04577_),
    .A3(_04578_),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04583_));
 sky130_fd_sc_hd__a22o_1 _11390_ (.A1(_04375_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_04582_),
    .B2(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__and2_1 _11391_ (.A(_04468_),
    .B(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _11392_ (.A(_04585_),
    .X(_00570_));
 sky130_fd_sc_hd__xnor2_1 _11393_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_04545_),
    .Y(_04586_));
 sky130_fd_sc_hd__a21oi_1 _11394_ (.A1(_04579_),
    .A2(_04582_),
    .B1(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__a31o_1 _11395_ (.A1(_04579_),
    .A2(_04582_),
    .A3(_04586_),
    .B1(_04396_),
    .X(_04588_));
 sky130_fd_sc_hd__o221a_1 _11396_ (.A1(_04431_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B1(_04587_),
    .B2(_04588_),
    .C1(_04539_),
    .X(_00571_));
 sky130_fd_sc_hd__and4b_1 _11397_ (.A_N(_04570_),
    .B(_04574_),
    .C(_04581_),
    .D(_04586_),
    .X(_04589_));
 sky130_fd_sc_hd__o41a_1 _11398_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A3(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A4(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_04565_),
    .X(_04590_));
 sky130_fd_sc_hd__or2_1 _11399_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04565_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04565_),
    .Y(_04592_));
 sky130_fd_sc_hd__and2_1 _11401_ (.A(_04591_),
    .B(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__o21ai_1 _11402_ (.A1(_04589_),
    .A2(_04590_),
    .B1(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__o31a_1 _11403_ (.A1(_04593_),
    .A2(_04589_),
    .A3(_04590_),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04595_));
 sky130_fd_sc_hd__a22o_1 _11404_ (.A1(_04375_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B1(_04594_),
    .B2(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__and2_1 _11405_ (.A(_04468_),
    .B(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _11406_ (.A(_04597_),
    .X(_00572_));
 sky130_fd_sc_hd__xnor2_1 _11407_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_04545_),
    .Y(_04598_));
 sky130_fd_sc_hd__a21oi_1 _11408_ (.A1(_04592_),
    .A2(_04594_),
    .B1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__a31o_1 _11409_ (.A1(_04592_),
    .A2(_04594_),
    .A3(_04598_),
    .B1(_04396_),
    .X(_04600_));
 sky130_fd_sc_hd__o221a_1 _11410_ (.A1(_04431_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B1(_04599_),
    .B2(_04600_),
    .C1(_04539_),
    .X(_00573_));
 sky130_fd_sc_hd__and2_1 _11411_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04601_));
 sky130_fd_sc_hd__nor2_1 _11412_ (.A(net282),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_2 _11413_ (.A1(_04601_),
    .A2(_04602_),
    .B1(_04391_),
    .Y(_04603_));
 sky130_fd_sc_hd__o211a_1 _11414_ (.A1(_04390_),
    .A2(net331),
    .B1(_04387_),
    .C1(_04603_),
    .X(_00574_));
 sky130_fd_sc_hd__and2b_1 _11415_ (.A_N(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04604_));
 sky130_fd_sc_hd__xnor2_1 _11416_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__xnor2_1 _11417_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__xor2_1 _11418_ (.A(_04601_),
    .B(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__or2_1 _11419_ (.A(_04444_),
    .B(net591),
    .X(_04608_));
 sky130_fd_sc_hd__o211a_1 _11420_ (.A1(_04442_),
    .A2(_04607_),
    .B1(_04608_),
    .C1(_04456_),
    .X(_00575_));
 sky130_fd_sc_hd__o21a_1 _11421_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_04412_),
    .X(_04609_));
 sky130_fd_sc_hd__xnor2_1 _11422_ (.A(net120),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__and2_1 _11423_ (.A(_04233_),
    .B(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__nor2_1 _11424_ (.A(_04233_),
    .B(_04610_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_1 _11425_ (.A(_04611_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__and2b_1 _11426_ (.A_N(_04605_),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_04614_));
 sky130_fd_sc_hd__a21o_1 _11427_ (.A1(_04601_),
    .A2(_04606_),
    .B1(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__nand2_1 _11428_ (.A(_04613_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__o21a_1 _11429_ (.A1(_04613_),
    .A2(_04615_),
    .B1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04617_));
 sky130_fd_sc_hd__a22o_1 _11430_ (.A1(_04375_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_04616_),
    .B2(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__and2_1 _11431_ (.A(_04468_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__clkbuf_1 _11432_ (.A(_04619_),
    .X(_00576_));
 sky130_fd_sc_hd__o31a_1 _11433_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A3(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_04412_),
    .X(_04620_));
 sky130_fd_sc_hd__xnor2_1 _11434_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__xnor2_1 _11435_ (.A(_04237_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__inv_2 _11436_ (.A(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__nand2_1 _11437_ (.A(_04233_),
    .B(_04610_),
    .Y(_04624_));
 sky130_fd_sc_hd__a21o_1 _11438_ (.A1(_04624_),
    .A2(_04615_),
    .B1(_04612_),
    .X(_04625_));
 sky130_fd_sc_hd__a21o_1 _11439_ (.A1(_04623_),
    .A2(_04625_),
    .B1(_04375_),
    .X(_04626_));
 sky130_fd_sc_hd__nor2_1 _11440_ (.A(_04623_),
    .B(_04625_),
    .Y(_04627_));
 sky130_fd_sc_hd__a2bb2o_1 _11441_ (.A1_N(_04626_),
    .A2_N(_04627_),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B2(_04375_),
    .X(_04628_));
 sky130_fd_sc_hd__and2_1 _11442_ (.A(_04468_),
    .B(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_04629_),
    .X(_00577_));
 sky130_fd_sc_hd__nor2_1 _11444_ (.A(_04237_),
    .B(_04621_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21oi_2 _11445_ (.A1(_04623_),
    .A2(_04625_),
    .B1(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__or4_4 _11446_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .C(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .D(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04632_));
 sky130_fd_sc_hd__nand2_1 _11447_ (.A(_04412_),
    .B(net652),
    .Y(_04633_));
 sky130_fd_sc_hd__xor2_2 _11448_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__xor2_2 _11449_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__xor2_1 _11450_ (.A(_04631_),
    .B(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__or2_1 _11451_ (.A(_04444_),
    .B(net513),
    .X(_04637_));
 sky130_fd_sc_hd__o211a_1 _11452_ (.A1(_04442_),
    .A2(_04636_),
    .B1(_04637_),
    .C1(_04456_),
    .X(_00578_));
 sky130_fd_sc_hd__o21a_1 _11453_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(net652),
    .B1(_04412_),
    .X(_04638_));
 sky130_fd_sc_hd__xor2_2 _11454_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__xnor2_1 _11455_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__inv_2 _11456_ (.A(_04634_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2_1 _11457_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__o21ai_1 _11458_ (.A1(_04631_),
    .A2(_04635_),
    .B1(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__xnor2_1 _11459_ (.A(_04640_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__or2_1 _11460_ (.A(_04444_),
    .B(net493),
    .X(_04645_));
 sky130_fd_sc_hd__o211a_1 _11461_ (.A1(_04442_),
    .A2(_04644_),
    .B1(_04645_),
    .C1(_04456_),
    .X(_00579_));
 sky130_fd_sc_hd__inv_2 _11462_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_04646_));
 sky130_fd_sc_hd__o31a_1 _11463_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A3(net652),
    .B1(_04413_),
    .X(_04647_));
 sky130_fd_sc_hd__xnor2_1 _11464_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__or2_1 _11465_ (.A(_04646_),
    .B(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__nand2_1 _11466_ (.A(_04646_),
    .B(_04648_),
    .Y(_04650_));
 sky130_fd_sc_hd__nand2_1 _11467_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__or2_1 _11468_ (.A(_04635_),
    .B(_04640_),
    .X(_04652_));
 sky130_fd_sc_hd__or2_1 _11469_ (.A(_04631_),
    .B(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__a22o_1 _11470_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .A2(_04641_),
    .B1(_04639_),
    .B2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_04654_));
 sky130_fd_sc_hd__o21ai_1 _11471_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(_04639_),
    .B1(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a31o_1 _11472_ (.A1(_04651_),
    .A2(_04653_),
    .A3(_04655_),
    .B1(_04374_),
    .X(_04656_));
 sky130_fd_sc_hd__a21oi_1 _11473_ (.A1(_04653_),
    .A2(_04655_),
    .B1(_04651_),
    .Y(_04657_));
 sky130_fd_sc_hd__a2bb2o_1 _11474_ (.A1_N(_04656_),
    .A2_N(_04657_),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B2(_04375_),
    .X(_04658_));
 sky130_fd_sc_hd__and2_1 _11475_ (.A(_04468_),
    .B(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__clkbuf_1 _11476_ (.A(_04659_),
    .X(_00580_));
 sky130_fd_sc_hd__inv_2 _11477_ (.A(_04649_),
    .Y(_04660_));
 sky130_fd_sc_hd__o41a_1 _11478_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A3(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A4(net652),
    .B1(_04412_),
    .X(_04661_));
 sky130_fd_sc_hd__xor2_1 _11479_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__nand2_1 _11480_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__nor2_1 _11481_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_04662_),
    .Y(_04664_));
 sky130_fd_sc_hd__inv_2 _11482_ (.A(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand2_1 _11483_ (.A(_04663_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__o21a_1 _11484_ (.A1(_04660_),
    .A2(_04657_),
    .B1(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__o31ai_1 _11485_ (.A1(_04660_),
    .A2(_04657_),
    .A3(_04666_),
    .B1(_04391_),
    .Y(_04668_));
 sky130_fd_sc_hd__o221a_1 _11486_ (.A1(_04431_),
    .A2(net406),
    .B1(_04667_),
    .B2(_04668_),
    .C1(_04539_),
    .X(_00581_));
 sky130_fd_sc_hd__inv_2 _11487_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_04669_));
 sky130_fd_sc_hd__or2_1 _11488_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_04670_));
 sky130_fd_sc_hd__or4_4 _11489_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .C(_04632_),
    .D(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__nand2_1 _11490_ (.A(_04413_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__xor2_1 _11491_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__nor2_1 _11492_ (.A(_04669_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__and2_1 _11493_ (.A(_04669_),
    .B(_04673_),
    .X(_04675_));
 sky130_fd_sc_hd__or2_2 _11494_ (.A(_04674_),
    .B(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__a21o_1 _11495_ (.A1(_04649_),
    .A2(_04663_),
    .B1(_04664_),
    .X(_04677_));
 sky130_fd_sc_hd__o31a_1 _11496_ (.A1(_04651_),
    .A2(_04655_),
    .A3(_04666_),
    .B1(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__or4_2 _11497_ (.A(_04631_),
    .B(_04651_),
    .C(_04652_),
    .D(_04666_),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _11498_ (.A(_04678_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xnor2_1 _11499_ (.A(_04676_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__or2_1 _11500_ (.A(_04444_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_04682_));
 sky130_fd_sc_hd__o211a_1 _11501_ (.A1(_04442_),
    .A2(_04681_),
    .B1(_04682_),
    .C1(_04456_),
    .X(_00582_));
 sky130_fd_sc_hd__o21a_1 _11502_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_04671_),
    .B1(_04413_),
    .X(_04683_));
 sky130_fd_sc_hd__xor2_2 _11503_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__xnor2_2 _11504_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _11505_ (.A(_04676_),
    .Y(_04686_));
 sky130_fd_sc_hd__a21o_1 _11506_ (.A1(_04686_),
    .A2(_04680_),
    .B1(_04674_),
    .X(_04687_));
 sky130_fd_sc_hd__nor2_1 _11507_ (.A(_04685_),
    .B(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21o_1 _11508_ (.A1(_04685_),
    .A2(_04687_),
    .B1(_04376_),
    .X(_04689_));
 sky130_fd_sc_hd__o221a_1 _11509_ (.A1(_04431_),
    .A2(net564),
    .B1(_04688_),
    .B2(_04689_),
    .C1(_04539_),
    .X(_00583_));
 sky130_fd_sc_hd__o31a_1 _11510_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A3(_04671_),
    .B1(_04412_),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_4 _11511_ (.A0(_04690_),
    .A1(_04061_),
    .S(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_04691_));
 sky130_fd_sc_hd__buf_6 _11512_ (.A(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__or4b_1 _11513_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(_04671_),
    .D_N(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_04693_));
 sky130_fd_sc_hd__or2b_4 _11514_ (.A(_04692_),
    .B_N(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__xnor2_4 _11515_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__nor2_1 _11516_ (.A(_04676_),
    .B(_04685_),
    .Y(_04696_));
 sky130_fd_sc_hd__a21o_1 _11517_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_04684_),
    .B1(_04674_),
    .X(_04697_));
 sky130_fd_sc_hd__o21ai_1 _11518_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_04684_),
    .B1(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__a21bo_1 _11519_ (.A1(_04680_),
    .A2(_04696_),
    .B1_N(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__or2b_1 _11520_ (.A(_04695_),
    .B_N(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__or2b_1 _11521_ (.A(_04699_),
    .B_N(_04695_),
    .X(_04701_));
 sky130_fd_sc_hd__and2_1 _11522_ (.A(_04375_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .X(_04702_));
 sky130_fd_sc_hd__a31o_1 _11523_ (.A1(_04378_),
    .A2(_04700_),
    .A3(_04701_),
    .B1(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__and2_1 _11524_ (.A(_04468_),
    .B(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_1 _11525_ (.A(_04704_),
    .X(_00584_));
 sky130_fd_sc_hd__nand2_1 _11526_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04692_),
    .Y(_04705_));
 sky130_fd_sc_hd__or2_1 _11527_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04692_),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_1 _11528_ (.A(_04705_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand2_1 _11529_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04694_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_1 _11530_ (.A(_04708_),
    .B(_04700_),
    .Y(_04709_));
 sky130_fd_sc_hd__nor2_1 _11531_ (.A(_04707_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__a21o_1 _11532_ (.A1(_04707_),
    .A2(_04709_),
    .B1(_04376_),
    .X(_04711_));
 sky130_fd_sc_hd__o221a_1 _11533_ (.A1(_04391_),
    .A2(net520),
    .B1(_04710_),
    .B2(_04711_),
    .C1(_04539_),
    .X(_00585_));
 sky130_fd_sc_hd__xnor2_1 _11534_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_04692_),
    .Y(_04712_));
 sky130_fd_sc_hd__nor2_1 _11535_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04692_),
    .Y(_04713_));
 sky130_fd_sc_hd__a21o_1 _11536_ (.A1(_04708_),
    .A2(_04705_),
    .B1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__or4_4 _11537_ (.A(_04676_),
    .B(_04685_),
    .C(_04695_),
    .D(_04707_),
    .X(_04715_));
 sky130_fd_sc_hd__a21o_1 _11538_ (.A1(_04678_),
    .A2(_04679_),
    .B1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__or3_1 _11539_ (.A(_04695_),
    .B(_04698_),
    .C(_04707_),
    .X(_04717_));
 sky130_fd_sc_hd__and3_1 _11540_ (.A(_04714_),
    .B(_04716_),
    .C(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _11541_ (.A(_04712_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__and2_1 _11542_ (.A(_04712_),
    .B(_04718_),
    .X(_04720_));
 sky130_fd_sc_hd__o21ai_1 _11543_ (.A1(_04719_),
    .A2(_04720_),
    .B1(_04391_),
    .Y(_04721_));
 sky130_fd_sc_hd__o211a_1 _11544_ (.A1(_04390_),
    .A2(net504),
    .B1(_04387_),
    .C1(_04721_),
    .X(_00586_));
 sky130_fd_sc_hd__xnor2_1 _11545_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_04692_),
    .Y(_04722_));
 sky130_fd_sc_hd__clkbuf_4 _11546_ (.A(_04692_),
    .X(_04723_));
 sky130_fd_sc_hd__a21o_1 _11547_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_04723_),
    .B1(_04719_),
    .X(_04724_));
 sky130_fd_sc_hd__xnor2_1 _11548_ (.A(_04722_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__or2_1 _11549_ (.A(_04378_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_04726_));
 sky130_fd_sc_hd__o211a_1 _11550_ (.A1(_04376_),
    .A2(_04725_),
    .B1(_04726_),
    .C1(_04456_),
    .X(_00587_));
 sky130_fd_sc_hd__and2_1 _11551_ (.A(_04396_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_04727_));
 sky130_fd_sc_hd__a31o_1 _11552_ (.A1(_04714_),
    .A2(_04716_),
    .A3(_04717_),
    .B1(_04712_),
    .X(_04728_));
 sky130_fd_sc_hd__o21bai_1 _11553_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(_04723_),
    .B1_N(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__o21ai_1 _11554_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_04723_),
    .Y(_04730_));
 sky130_fd_sc_hd__xnor2_1 _11555_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_04723_),
    .Y(_04731_));
 sky130_fd_sc_hd__a21oi_1 _11556_ (.A1(_04729_),
    .A2(_04730_),
    .B1(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__a31o_1 _11557_ (.A1(_04731_),
    .A2(_04729_),
    .A3(_04730_),
    .B1(_04396_),
    .X(_04733_));
 sky130_fd_sc_hd__nor2_1 _11558_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__o21a_1 _11559_ (.A1(_04727_),
    .A2(_04734_),
    .B1(_02132_),
    .X(_00588_));
 sky130_fd_sc_hd__xnor2_1 _11560_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_04723_),
    .Y(_04735_));
 sky130_fd_sc_hd__a21o_1 _11561_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_04723_),
    .B1(_04732_),
    .X(_04736_));
 sky130_fd_sc_hd__xnor2_1 _11562_ (.A(_04735_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__or2_1 _11563_ (.A(_04378_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(_04738_));
 sky130_fd_sc_hd__clkbuf_4 _11564_ (.A(_04455_),
    .X(_04739_));
 sky130_fd_sc_hd__o211a_1 _11565_ (.A1(_04376_),
    .A2(_04737_),
    .B1(_04738_),
    .C1(_04739_),
    .X(_00589_));
 sky130_fd_sc_hd__or2_1 _11566_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04723_),
    .X(_04740_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04723_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand2_1 _11568_ (.A(_04740_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__or4_1 _11569_ (.A(_04728_),
    .B(_04722_),
    .C(_04731_),
    .D(_04735_),
    .X(_04743_));
 sky130_fd_sc_hd__o21ai_1 _11570_ (.A1(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_04723_),
    .Y(_04744_));
 sky130_fd_sc_hd__and3_1 _11571_ (.A(_04730_),
    .B(_04743_),
    .C(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__xor2_1 _11572_ (.A(_04742_),
    .B(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A1(_04746_),
    .S(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04747_));
 sky130_fd_sc_hd__and2_4 _11574_ (.A(_04468_),
    .B(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _11575_ (.A(_04748_),
    .X(_00590_));
 sky130_fd_sc_hd__o21ai_1 _11576_ (.A1(_04742_),
    .A2(_04745_),
    .B1(_04741_),
    .Y(_04749_));
 sky130_fd_sc_hd__xnor2_1 _11577_ (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_04723_),
    .Y(_04750_));
 sky130_fd_sc_hd__xnor2_1 _11578_ (.A(_04749_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__or2_1 _11579_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_04378_),
    .X(_04752_));
 sky130_fd_sc_hd__o211a_1 _11580_ (.A1(_04376_),
    .A2(_04751_),
    .B1(_04752_),
    .C1(_04739_),
    .X(_00591_));
 sky130_fd_sc_hd__and2_1 _11581_ (.A(_04391_),
    .B(_02310_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_1 _11582_ (.A(_04753_),
    .X(_00592_));
 sky130_fd_sc_hd__inv_2 _11583_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_04754_));
 sky130_fd_sc_hd__clkbuf_4 _11584_ (.A(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__clkbuf_4 _11585_ (.A(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__clkbuf_4 _11586_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_04757_));
 sky130_fd_sc_hd__clkbuf_4 _11587_ (.A(_04757_),
    .X(_04758_));
 sky130_fd_sc_hd__or2_1 _11588_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__o211a_1 _11589_ (.A1(_04756_),
    .A2(net143),
    .B1(_04387_),
    .C1(_04759_),
    .X(_00593_));
 sky130_fd_sc_hd__or2_1 _11590_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_04758_),
    .X(_04760_));
 sky130_fd_sc_hd__o211a_1 _11591_ (.A1(_04756_),
    .A2(net128),
    .B1(_04387_),
    .C1(_04760_),
    .X(_00594_));
 sky130_fd_sc_hd__or2_1 _11592_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B(_04758_),
    .X(_04761_));
 sky130_fd_sc_hd__o211a_1 _11593_ (.A1(_04756_),
    .A2(net122),
    .B1(_04387_),
    .C1(_04761_),
    .X(_00595_));
 sky130_fd_sc_hd__clkbuf_4 _11594_ (.A(_03619_),
    .X(_04762_));
 sky130_fd_sc_hd__or2_1 _11595_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(_04758_),
    .X(_04763_));
 sky130_fd_sc_hd__o211a_1 _11596_ (.A1(_04756_),
    .A2(net151),
    .B1(_04762_),
    .C1(_04763_),
    .X(_00596_));
 sky130_fd_sc_hd__or2_1 _11597_ (.A(net162),
    .B(_04758_),
    .X(_04764_));
 sky130_fd_sc_hd__o211a_1 _11598_ (.A1(_04756_),
    .A2(net166),
    .B1(_04762_),
    .C1(_04764_),
    .X(_00597_));
 sky130_fd_sc_hd__buf_2 _11599_ (.A(_04757_),
    .X(_04765_));
 sky130_fd_sc_hd__or2_1 _11600_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__o211a_1 _11601_ (.A1(_04756_),
    .A2(net134),
    .B1(_04762_),
    .C1(_04766_),
    .X(_00598_));
 sky130_fd_sc_hd__or2_1 _11602_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_04765_),
    .X(_04767_));
 sky130_fd_sc_hd__o211a_1 _11603_ (.A1(_04756_),
    .A2(net138),
    .B1(_04762_),
    .C1(_04767_),
    .X(_00599_));
 sky130_fd_sc_hd__or2_1 _11604_ (.A(_04758_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(_04768_));
 sky130_fd_sc_hd__o211a_1 _11605_ (.A1(_04756_),
    .A2(net161),
    .B1(_04762_),
    .C1(_04768_),
    .X(_00600_));
 sky130_fd_sc_hd__clkbuf_4 _11606_ (.A(_04765_),
    .X(_04769_));
 sky130_fd_sc_hd__buf_2 _11607_ (.A(_04757_),
    .X(_04770_));
 sky130_fd_sc_hd__clkbuf_4 _11608_ (.A(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__nand2_1 _11609_ (.A(_04771_),
    .B(net274),
    .Y(_04772_));
 sky130_fd_sc_hd__o211a_1 _11610_ (.A1(_04769_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B1(_04762_),
    .C1(_04772_),
    .X(_00601_));
 sky130_fd_sc_hd__clkbuf_4 _11611_ (.A(_04770_),
    .X(_04773_));
 sky130_fd_sc_hd__nand2_1 _11612_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .Y(_04774_));
 sky130_fd_sc_hd__or2_1 _11613_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(_04775_));
 sky130_fd_sc_hd__a21oi_1 _11614_ (.A1(_04774_),
    .A2(_04775_),
    .B1(_04445_),
    .Y(_04776_));
 sky130_fd_sc_hd__a31o_1 _11615_ (.A1(_04445_),
    .A2(_04774_),
    .A3(_04775_),
    .B1(_04755_),
    .X(_04777_));
 sky130_fd_sc_hd__o221a_1 _11616_ (.A1(_04773_),
    .A2(net509),
    .B1(_04776_),
    .B2(_04777_),
    .C1(_04539_),
    .X(_00602_));
 sky130_fd_sc_hd__and3_1 _11617_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(_04778_));
 sky130_fd_sc_hd__a21oi_1 _11618_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .Y(_04779_));
 sky130_fd_sc_hd__or2_1 _11619_ (.A(_04778_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_1 _11620_ (.A(_04776_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__a21o_1 _11621_ (.A1(_04776_),
    .A2(_04780_),
    .B1(_04755_),
    .X(_04782_));
 sky130_fd_sc_hd__o221a_1 _11622_ (.A1(_04773_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B1(_04781_),
    .B2(_04782_),
    .C1(_04539_),
    .X(_00603_));
 sky130_fd_sc_hd__nand2_1 _11623_ (.A(_04445_),
    .B(_04778_),
    .Y(_04783_));
 sky130_fd_sc_hd__o31a_1 _11624_ (.A1(_04445_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A3(_04775_),
    .B1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__and2_1 _11625_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_4 _11626_ (.A(_04770_),
    .X(_04786_));
 sky130_fd_sc_hd__o21ai_1 _11627_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_04784_),
    .B1(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__clkbuf_4 _11628_ (.A(_04538_),
    .X(_04788_));
 sky130_fd_sc_hd__o221a_1 _11629_ (.A1(_04773_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_04785_),
    .B2(_04787_),
    .C1(_04788_),
    .X(_00604_));
 sky130_fd_sc_hd__or3_1 _11630_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(_04775_),
    .X(_04789_));
 sky130_fd_sc_hd__nand2_1 _11631_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_04778_),
    .Y(_04790_));
 sky130_fd_sc_hd__mux2_1 _11632_ (.A0(_04789_),
    .A1(_04790_),
    .S(_04445_),
    .X(_04791_));
 sky130_fd_sc_hd__and2_1 _11633_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__o21ai_1 _11634_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_04791_),
    .B1(_04786_),
    .Y(_04793_));
 sky130_fd_sc_hd__o221a_1 _11635_ (.A1(_04773_),
    .A2(net476),
    .B1(_04792_),
    .B2(_04793_),
    .C1(_04788_),
    .X(_00605_));
 sky130_fd_sc_hd__inv_2 _11636_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_04794_));
 sky130_fd_sc_hd__clkbuf_4 _11637_ (.A(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__o21ai_1 _11638_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_04789_),
    .B1(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__a31o_1 _11639_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A3(_04778_),
    .B1(_04795_),
    .X(_04797_));
 sky130_fd_sc_hd__inv_2 _11640_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .Y(_04798_));
 sky130_fd_sc_hd__a21oi_1 _11641_ (.A1(_04796_),
    .A2(_04797_),
    .B1(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__a31o_1 _11642_ (.A1(_04798_),
    .A2(_04796_),
    .A3(_04797_),
    .B1(_04755_),
    .X(_04800_));
 sky130_fd_sc_hd__o221a_1 _11643_ (.A1(_04773_),
    .A2(net625),
    .B1(_04799_),
    .B2(_04800_),
    .C1(_04788_),
    .X(_00606_));
 sky130_fd_sc_hd__and4_1 _11644_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .D(_04778_),
    .X(_04801_));
 sky130_fd_sc_hd__or3_1 _11645_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_04789_),
    .X(_04802_));
 sky130_fd_sc_hd__inv_2 _11646_ (.A(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(_04801_),
    .A1(_04803_),
    .S(_04795_),
    .X(_04804_));
 sky130_fd_sc_hd__xnor2_1 _11648_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand2_1 _11649_ (.A(_04771_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__o211a_1 _11650_ (.A1(_04769_),
    .A2(net560),
    .B1(_04762_),
    .C1(_04806_),
    .X(_00607_));
 sky130_fd_sc_hd__or2_1 _11651_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_04802_),
    .X(_04807_));
 sky130_fd_sc_hd__and2_1 _11652_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_04801_),
    .X(_04808_));
 sky130_fd_sc_hd__nand2_1 _11653_ (.A(_04445_),
    .B(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__o21a_1 _11654_ (.A1(_04445_),
    .A2(_04807_),
    .B1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__o21ai_1 _11655_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_04810_),
    .B1(_04770_),
    .Y(_04811_));
 sky130_fd_sc_hd__a21o_1 _11656_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_04810_),
    .B1(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__o211a_1 _11657_ (.A1(_04769_),
    .A2(net572),
    .B1(_04762_),
    .C1(_04812_),
    .X(_00608_));
 sky130_fd_sc_hd__nand3_1 _11658_ (.A(_04445_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_04808_),
    .Y(_04813_));
 sky130_fd_sc_hd__o31a_1 _11659_ (.A1(_04445_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A3(_04807_),
    .B1(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__and2_1 _11660_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__o21ai_1 _11661_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_04814_),
    .B1(_04786_),
    .Y(_04816_));
 sky130_fd_sc_hd__o221a_1 _11662_ (.A1(_04773_),
    .A2(net566),
    .B1(_04815_),
    .B2(_04816_),
    .C1(_04788_),
    .X(_00609_));
 sky130_fd_sc_hd__and3_1 _11663_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_04808_),
    .X(_04817_));
 sky130_fd_sc_hd__inv_2 _11664_ (.A(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__or3_1 _11665_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_04807_),
    .X(_04819_));
 sky130_fd_sc_hd__mux2_1 _11666_ (.A0(_04818_),
    .A1(_04819_),
    .S(_04795_),
    .X(_04820_));
 sky130_fd_sc_hd__nor2_1 _11667_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21o_1 _11668_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_04820_),
    .B1(_04755_),
    .X(_04822_));
 sky130_fd_sc_hd__o221a_1 _11669_ (.A1(_04773_),
    .A2(net606),
    .B1(_04821_),
    .B2(_04822_),
    .C1(_04788_),
    .X(_00610_));
 sky130_fd_sc_hd__o21a_1 _11670_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_04819_),
    .B1(_04795_),
    .X(_04823_));
 sky130_fd_sc_hd__a21o_1 _11671_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_04817_),
    .B1(_04795_),
    .X(_04824_));
 sky130_fd_sc_hd__or2b_1 _11672_ (.A(_04823_),
    .B_N(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__nor2_1 _11673_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__a21o_1 _11674_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_04825_),
    .B1(_04755_),
    .X(_04827_));
 sky130_fd_sc_hd__o221a_1 _11675_ (.A1(_04773_),
    .A2(net522),
    .B1(_04826_),
    .B2(_04827_),
    .C1(_04788_),
    .X(_00611_));
 sky130_fd_sc_hd__a21oi_1 _11676_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_04824_),
    .B1(_04823_),
    .Y(_04828_));
 sky130_fd_sc_hd__buf_2 _11677_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_04829_));
 sky130_fd_sc_hd__or2_1 _11678_ (.A(_04765_),
    .B(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__o211a_1 _11679_ (.A1(_04756_),
    .A2(_04828_),
    .B1(_04830_),
    .C1(_04739_),
    .X(_00612_));
 sky130_fd_sc_hd__inv_2 _11680_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .Y(_04831_));
 sky130_fd_sc_hd__nor2_1 _11681_ (.A(_04831_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_04832_));
 sky130_fd_sc_hd__a21o_1 _11682_ (.A1(_04831_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_04755_),
    .X(_04833_));
 sky130_fd_sc_hd__o221a_1 _11683_ (.A1(_04773_),
    .A2(net391),
    .B1(_04832_),
    .B2(_04833_),
    .C1(_04788_),
    .X(_00613_));
 sky130_fd_sc_hd__and2b_1 _11684_ (.A_N(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_04834_));
 sky130_fd_sc_hd__xnor2_1 _11685_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__xnor2_1 _11686_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__xor2_1 _11687_ (.A(_04832_),
    .B(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _11688_ (.A(_04765_),
    .B(net633),
    .X(_04838_));
 sky130_fd_sc_hd__o211a_1 _11689_ (.A1(_04756_),
    .A2(_04837_),
    .B1(_04838_),
    .C1(_04739_),
    .X(_00614_));
 sky130_fd_sc_hd__and2_1 _11690_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_04835_),
    .X(_04839_));
 sky130_fd_sc_hd__nor2_1 _11691_ (.A(_04832_),
    .B(_04836_),
    .Y(_04840_));
 sky130_fd_sc_hd__o21ba_1 _11692_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1_N(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_04841_));
 sky130_fd_sc_hd__xnor2_1 _11693_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__or2_1 _11694_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__nand2_1 _11695_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_04842_),
    .Y(_04844_));
 sky130_fd_sc_hd__and2_1 _11696_ (.A(_04843_),
    .B(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__o21ai_1 _11697_ (.A1(_04839_),
    .A2(_04840_),
    .B1(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__o31a_1 _11698_ (.A1(_04839_),
    .A2(_04840_),
    .A3(_04845_),
    .B1(_04757_),
    .X(_04847_));
 sky130_fd_sc_hd__a22oi_1 _11699_ (.A1(_04754_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_04846_),
    .B2(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__and2b_1 _11700_ (.A_N(_04848_),
    .B(_03118_),
    .X(_04849_));
 sky130_fd_sc_hd__clkbuf_1 _11701_ (.A(_04849_),
    .X(_00615_));
 sky130_fd_sc_hd__buf_2 _11702_ (.A(_01252_),
    .X(_04850_));
 sky130_fd_sc_hd__o31a_1 _11703_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A3(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_04794_),
    .X(_04851_));
 sky130_fd_sc_hd__xnor2_1 _11704_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__and2_1 _11705_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__nor2_1 _11706_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_04852_),
    .Y(_04854_));
 sky130_fd_sc_hd__nor2_1 _11707_ (.A(_04853_),
    .B(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__a21boi_1 _11708_ (.A1(_04844_),
    .A2(_04846_),
    .B1_N(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_1 _11709_ (.A(_04754_),
    .B(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _11710_ (.A(_04844_),
    .B(_04846_),
    .Y(_04858_));
 sky130_fd_sc_hd__nor2_1 _11711_ (.A(_04855_),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__a2bb2o_1 _11712_ (.A1_N(_04857_),
    .A2_N(_04859_),
    .B1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B2(_04754_),
    .X(_04860_));
 sky130_fd_sc_hd__and2_1 _11713_ (.A(_04850_),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_1 _11714_ (.A(_04861_),
    .X(_00616_));
 sky130_fd_sc_hd__clkbuf_4 _11715_ (.A(_04754_),
    .X(_04862_));
 sky130_fd_sc_hd__or2_1 _11716_ (.A(_04853_),
    .B(_04856_),
    .X(_04863_));
 sky130_fd_sc_hd__or4_2 _11717_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .D(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_04864_));
 sky130_fd_sc_hd__a21oi_1 _11718_ (.A1(_04794_),
    .A2(_04864_),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .Y(_04865_));
 sky130_fd_sc_hd__and3_1 _11719_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_04794_),
    .C(_04864_),
    .X(_04866_));
 sky130_fd_sc_hd__or2_1 _11720_ (.A(_04865_),
    .B(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__and2_1 _11721_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__nor2_1 _11722_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_04867_),
    .Y(_04869_));
 sky130_fd_sc_hd__nor2_1 _11723_ (.A(_04868_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__xor2_1 _11724_ (.A(_04863_),
    .B(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__or2_1 _11725_ (.A(_04765_),
    .B(net497),
    .X(_04872_));
 sky130_fd_sc_hd__o211a_1 _11726_ (.A1(_04862_),
    .A2(_04871_),
    .B1(_04872_),
    .C1(_04739_),
    .X(_00617_));
 sky130_fd_sc_hd__o21a_1 _11727_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(_04864_),
    .B1(_04794_),
    .X(_04873_));
 sky130_fd_sc_hd__xor2_1 _11728_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__and2b_1 _11729_ (.A_N(_04874_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_04875_));
 sky130_fd_sc_hd__or2b_1 _11730_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B_N(_04874_),
    .X(_04876_));
 sky130_fd_sc_hd__and2b_1 _11731_ (.A_N(_04875_),
    .B(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__a21oi_1 _11732_ (.A1(_04863_),
    .A2(_04870_),
    .B1(_04868_),
    .Y(_04878_));
 sky130_fd_sc_hd__xnor2_1 _11733_ (.A(_04877_),
    .B(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_1 _11734_ (.A(_04765_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_04880_));
 sky130_fd_sc_hd__o211a_1 _11735_ (.A1(_04862_),
    .A2(_04879_),
    .B1(_04880_),
    .C1(_04739_),
    .X(_00618_));
 sky130_fd_sc_hd__and2_1 _11736_ (.A(_04870_),
    .B(_04877_),
    .X(_04881_));
 sky130_fd_sc_hd__and2_1 _11737_ (.A(_04863_),
    .B(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__o21a_1 _11738_ (.A1(_04868_),
    .A2(_04875_),
    .B1(_04876_),
    .X(_04883_));
 sky130_fd_sc_hd__o31a_1 _11739_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A3(_04864_),
    .B1(_04794_),
    .X(_04884_));
 sky130_fd_sc_hd__xnor2_1 _11740_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _11741_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__or2_1 _11742_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_04885_),
    .X(_04887_));
 sky130_fd_sc_hd__and2_1 _11743_ (.A(_04886_),
    .B(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__o21ai_1 _11744_ (.A1(_04882_),
    .A2(_04883_),
    .B1(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__o31a_1 _11745_ (.A1(_04888_),
    .A2(_04882_),
    .A3(_04883_),
    .B1(_04757_),
    .X(_04890_));
 sky130_fd_sc_hd__a22o_1 _11746_ (.A1(_04754_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_04889_),
    .B2(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__and2_1 _11747_ (.A(_04850_),
    .B(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__clkbuf_1 _11748_ (.A(_04892_),
    .X(_00619_));
 sky130_fd_sc_hd__a21o_1 _11749_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_04794_),
    .B1(_04884_),
    .X(_04893_));
 sky130_fd_sc_hd__xor2_1 _11750_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__or2b_1 _11751_ (.A(_04894_),
    .B_N(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_04895_));
 sky130_fd_sc_hd__or2b_1 _11752_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B_N(_04894_),
    .X(_04896_));
 sky130_fd_sc_hd__and2_1 _11753_ (.A(_04895_),
    .B(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__a21oi_1 _11754_ (.A1(_04886_),
    .A2(_04889_),
    .B1(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__a31o_1 _11755_ (.A1(_04886_),
    .A2(_04889_),
    .A3(_04897_),
    .B1(_04755_),
    .X(_04899_));
 sky130_fd_sc_hd__o221a_1 _11756_ (.A1(_04773_),
    .A2(net443),
    .B1(_04898_),
    .B2(_04899_),
    .C1(_04788_),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _11757_ (.A(_04886_),
    .B(_04895_),
    .Y(_04900_));
 sky130_fd_sc_hd__a32o_1 _11758_ (.A1(_04888_),
    .A2(_04883_),
    .A3(_04897_),
    .B1(_04900_),
    .B2(_04896_),
    .X(_04901_));
 sky130_fd_sc_hd__o2111a_1 _11759_ (.A1(_04853_),
    .A2(_04856_),
    .B1(_04888_),
    .C1(_04881_),
    .D1(_04897_),
    .X(_04902_));
 sky130_fd_sc_hd__or4_1 _11760_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .D(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_04903_));
 sky130_fd_sc_hd__or2_1 _11761_ (.A(_04864_),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(_04795_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__xor2_1 _11763_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_1 _11764_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__or2_1 _11765_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_04906_),
    .X(_04908_));
 sky130_fd_sc_hd__and2_1 _11766_ (.A(_04907_),
    .B(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__o21ai_2 _11767_ (.A1(_04901_),
    .A2(_04902_),
    .B1(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__or3_1 _11768_ (.A(_04909_),
    .B(_04901_),
    .C(_04902_),
    .X(_04911_));
 sky130_fd_sc_hd__a21o_1 _11769_ (.A1(_04910_),
    .A2(_04911_),
    .B1(_04862_),
    .X(_04912_));
 sky130_fd_sc_hd__o211a_1 _11770_ (.A1(_04769_),
    .A2(net389),
    .B1(_04762_),
    .C1(_04912_),
    .X(_00621_));
 sky130_fd_sc_hd__o21ai_1 _11771_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_04904_),
    .B1(_04794_),
    .Y(_04913_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(_04913_),
    .A1(_04795_),
    .S(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_04914_));
 sky130_fd_sc_hd__buf_2 _11773_ (.A(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__or3b_1 _11774_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_04904_),
    .C_N(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_04916_));
 sky130_fd_sc_hd__a21o_1 _11775_ (.A1(_04915_),
    .A2(_04916_),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_04917_));
 sky130_fd_sc_hd__nand3_1 _11776_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_04915_),
    .C(_04916_),
    .Y(_04918_));
 sky130_fd_sc_hd__nand2_1 _11777_ (.A(_04917_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__and3_1 _11778_ (.A(_04907_),
    .B(_04910_),
    .C(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__a21oi_1 _11779_ (.A1(_04907_),
    .A2(_04910_),
    .B1(_04919_),
    .Y(_04921_));
 sky130_fd_sc_hd__o21ai_1 _11780_ (.A1(_04920_),
    .A2(_04921_),
    .B1(_04771_),
    .Y(_04922_));
 sky130_fd_sc_hd__o211a_1 _11781_ (.A1(_04769_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_04762_),
    .C1(_04922_),
    .X(_00622_));
 sky130_fd_sc_hd__nand2_1 _11782_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04915_),
    .Y(_04923_));
 sky130_fd_sc_hd__or2_1 _11783_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04915_),
    .X(_04924_));
 sky130_fd_sc_hd__nand2_1 _11784_ (.A(_04923_),
    .B(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__inv_2 _11785_ (.A(_04917_),
    .Y(_04926_));
 sky130_fd_sc_hd__a31o_1 _11786_ (.A1(_04907_),
    .A2(_04910_),
    .A3(_04918_),
    .B1(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__xor2_1 _11787_ (.A(_04925_),
    .B(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__or2_1 _11788_ (.A(_04765_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_04929_));
 sky130_fd_sc_hd__o211a_1 _11789_ (.A1(_04862_),
    .A2(_04928_),
    .B1(_04929_),
    .C1(_04739_),
    .X(_00623_));
 sky130_fd_sc_hd__clkbuf_4 _11790_ (.A(_04915_),
    .X(_04930_));
 sky130_fd_sc_hd__xor2_1 _11791_ (.A(_04557_),
    .B(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__o21a_1 _11792_ (.A1(_04925_),
    .A2(_04927_),
    .B1(_04923_),
    .X(_04932_));
 sky130_fd_sc_hd__and2_1 _11793_ (.A(_04931_),
    .B(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__o21ai_1 _11794_ (.A1(_04931_),
    .A2(_04932_),
    .B1(_04786_),
    .Y(_04934_));
 sky130_fd_sc_hd__o221a_1 _11795_ (.A1(_04771_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_04933_),
    .B2(_04934_),
    .C1(_04788_),
    .X(_00624_));
 sky130_fd_sc_hd__o21ai_1 _11796_ (.A1(_04557_),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_04915_),
    .Y(_04935_));
 sky130_fd_sc_hd__xnor2_1 _11797_ (.A(_04557_),
    .B(_04915_),
    .Y(_04936_));
 sky130_fd_sc_hd__a2111o_1 _11798_ (.A1(_04907_),
    .A2(_04918_),
    .B1(_04925_),
    .C1(_04936_),
    .D1(_04926_),
    .X(_04937_));
 sky130_fd_sc_hd__and2_1 _11799_ (.A(_04917_),
    .B(_04918_),
    .X(_04938_));
 sky130_fd_sc_hd__nor2_1 _11800_ (.A(_04925_),
    .B(_04936_),
    .Y(_04939_));
 sky130_fd_sc_hd__o2111ai_1 _11801_ (.A1(_04901_),
    .A2(_04902_),
    .B1(_04938_),
    .C1(_04939_),
    .D1(_04909_),
    .Y(_04940_));
 sky130_fd_sc_hd__and3_1 _11802_ (.A(_04935_),
    .B(_04937_),
    .C(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_1 _11803_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04930_),
    .Y(_04942_));
 sky130_fd_sc_hd__and2_1 _11804_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_04915_),
    .X(_04943_));
 sky130_fd_sc_hd__or2_1 _11805_ (.A(_04942_),
    .B(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__xor2_1 _11806_ (.A(_04941_),
    .B(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__or2_1 _11807_ (.A(_04765_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_04946_));
 sky130_fd_sc_hd__o211a_1 _11808_ (.A1(_04862_),
    .A2(_04945_),
    .B1(_04946_),
    .C1(_04739_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_1 _11809_ (.A(_04941_),
    .B(_04944_),
    .Y(_04947_));
 sky130_fd_sc_hd__xnor2_1 _11810_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_04930_),
    .Y(_04948_));
 sky130_fd_sc_hd__o21a_1 _11811_ (.A1(_04943_),
    .A2(_04947_),
    .B1(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__o31ai_1 _11812_ (.A1(_04943_),
    .A2(_04947_),
    .A3(_04948_),
    .B1(_04758_),
    .Y(_04950_));
 sky130_fd_sc_hd__o221a_1 _11813_ (.A1(_04771_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_04949_),
    .B2(_04950_),
    .C1(_04788_),
    .X(_00626_));
 sky130_fd_sc_hd__and2_1 _11814_ (.A(_04755_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .X(_04951_));
 sky130_fd_sc_hd__nor2_1 _11815_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .Y(_04952_));
 sky130_fd_sc_hd__or2b_1 _11816_ (.A(_04952_),
    .B_N(_04930_),
    .X(_04953_));
 sky130_fd_sc_hd__or3_1 _11817_ (.A(_04941_),
    .B(_04944_),
    .C(_04948_),
    .X(_04954_));
 sky130_fd_sc_hd__nor2_1 _11818_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04930_),
    .Y(_04955_));
 sky130_fd_sc_hd__and2_1 _11819_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_04915_),
    .X(_04956_));
 sky130_fd_sc_hd__or2_1 _11820_ (.A(_04955_),
    .B(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__a21oi_1 _11821_ (.A1(_04953_),
    .A2(_04954_),
    .B1(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__a31o_1 _11822_ (.A1(_04957_),
    .A2(_04953_),
    .A3(_04954_),
    .B1(_04754_),
    .X(_04959_));
 sky130_fd_sc_hd__nor2_1 _11823_ (.A(_04958_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__buf_6 _11824_ (.A(_01794_),
    .X(_04961_));
 sky130_fd_sc_hd__o21a_1 _11825_ (.A1(_04951_),
    .A2(_04960_),
    .B1(_04961_),
    .X(_00627_));
 sky130_fd_sc_hd__xnor2_1 _11826_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_04930_),
    .Y(_04962_));
 sky130_fd_sc_hd__o21a_1 _11827_ (.A1(_04956_),
    .A2(_04958_),
    .B1(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__o31ai_1 _11828_ (.A1(_04956_),
    .A2(_04958_),
    .A3(_04962_),
    .B1(_04758_),
    .Y(_04964_));
 sky130_fd_sc_hd__clkbuf_4 _11829_ (.A(_04538_),
    .X(_04965_));
 sky130_fd_sc_hd__o221a_1 _11830_ (.A1(_04771_),
    .A2(net589),
    .B1(_04963_),
    .B2(_04964_),
    .C1(_04965_),
    .X(_00628_));
 sky130_fd_sc_hd__or2_1 _11831_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04930_),
    .X(_04966_));
 sky130_fd_sc_hd__nand2_1 _11832_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_04930_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand2_1 _11833_ (.A(_04966_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_1 _11834_ (.A(_04957_),
    .B(_04962_),
    .X(_04969_));
 sky130_fd_sc_hd__or4_1 _11835_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .D(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_04970_));
 sky130_fd_sc_hd__a2bb2o_1 _11836_ (.A1_N(_04954_),
    .A2_N(_04969_),
    .B1(_04970_),
    .B2(_04930_),
    .X(_04971_));
 sky130_fd_sc_hd__xnor2_1 _11837_ (.A(_04968_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A1(_04972_),
    .S(_04757_),
    .X(_04973_));
 sky130_fd_sc_hd__and2_1 _11839_ (.A(_04850_),
    .B(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__clkbuf_1 _11840_ (.A(_04974_),
    .X(_00629_));
 sky130_fd_sc_hd__a21boi_1 _11841_ (.A1(_04966_),
    .A2(_04971_),
    .B1_N(_04967_),
    .Y(_04975_));
 sky130_fd_sc_hd__xnor2_1 _11842_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_04930_),
    .Y(_04976_));
 sky130_fd_sc_hd__xnor2_1 _11843_ (.A(_04975_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__o21ai_1 _11844_ (.A1(_04786_),
    .A2(net414),
    .B1(_01794_),
    .Y(_04978_));
 sky130_fd_sc_hd__a21oi_1 _11845_ (.A1(_04769_),
    .A2(_04977_),
    .B1(_04978_),
    .Y(_00630_));
 sky130_fd_sc_hd__clkbuf_4 _11846_ (.A(_03619_),
    .X(_04979_));
 sky130_fd_sc_hd__and2_1 _11847_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_04980_));
 sky130_fd_sc_hd__nor2_1 _11848_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .Y(_04981_));
 sky130_fd_sc_hd__o21ai_1 _11849_ (.A1(_04980_),
    .A2(_04981_),
    .B1(_04786_),
    .Y(_04982_));
 sky130_fd_sc_hd__o211a_1 _11850_ (.A1(_04769_),
    .A2(net271),
    .B1(_04979_),
    .C1(_04982_),
    .X(_00631_));
 sky130_fd_sc_hd__and2b_1 _11851_ (.A_N(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_04983_));
 sky130_fd_sc_hd__xnor2_1 _11852_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__xnor2_1 _11853_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__nor2_1 _11854_ (.A(_04980_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__and2_1 _11855_ (.A(_04980_),
    .B(_04985_),
    .X(_04987_));
 sky130_fd_sc_hd__o21ai_1 _11856_ (.A1(_04986_),
    .A2(_04987_),
    .B1(_04786_),
    .Y(_04988_));
 sky130_fd_sc_hd__o211a_1 _11857_ (.A1(_04769_),
    .A2(net312),
    .B1(_04979_),
    .C1(_04988_),
    .X(_00632_));
 sky130_fd_sc_hd__and2b_1 _11858_ (.A_N(_04984_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_04989_));
 sky130_fd_sc_hd__inv_2 _11859_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_04990_));
 sky130_fd_sc_hd__o21a_1 _11860_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_04794_),
    .X(_04991_));
 sky130_fd_sc_hd__xnor2_1 _11861_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__xnor2_1 _11862_ (.A(_04990_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__o21bai_2 _11863_ (.A1(_04989_),
    .A2(_04987_),
    .B1_N(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__or3b_1 _11864_ (.A(_04989_),
    .B(_04987_),
    .C_N(_04993_),
    .X(_04995_));
 sky130_fd_sc_hd__inv_2 _11865_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_04996_));
 sky130_fd_sc_hd__nor2_1 _11866_ (.A(_04757_),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__a31o_1 _11867_ (.A1(_04770_),
    .A2(_04994_),
    .A3(_04995_),
    .B1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__and2_1 _11868_ (.A(_04850_),
    .B(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__clkbuf_1 _11869_ (.A(_04999_),
    .X(_00633_));
 sky130_fd_sc_hd__inv_2 _11870_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_05000_));
 sky130_fd_sc_hd__or2_1 _11871_ (.A(_04990_),
    .B(_04992_),
    .X(_05001_));
 sky130_fd_sc_hd__inv_2 _11872_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_05002_));
 sky130_fd_sc_hd__o31a_1 _11873_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A3(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_04794_),
    .X(_05003_));
 sky130_fd_sc_hd__xnor2_1 _11874_ (.A(_04557_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(_05002_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__and2_1 _11876_ (.A(_05002_),
    .B(_05004_),
    .X(_05006_));
 sky130_fd_sc_hd__or2_1 _11877_ (.A(_05005_),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__and3_1 _11878_ (.A(_05001_),
    .B(_04994_),
    .C(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__a21oi_1 _11879_ (.A1(_05001_),
    .A2(_04994_),
    .B1(_05007_),
    .Y(_05009_));
 sky130_fd_sc_hd__or3_1 _11880_ (.A(_04754_),
    .B(_05008_),
    .C(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__o21a_1 _11881_ (.A1(_04770_),
    .A2(_05000_),
    .B1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__and2b_1 _11882_ (.A_N(_05011_),
    .B(_03118_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(_05012_),
    .X(_00634_));
 sky130_fd_sc_hd__nor2_1 _11884_ (.A(_05005_),
    .B(_05009_),
    .Y(_05013_));
 sky130_fd_sc_hd__inv_2 _11885_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_05014_));
 sky130_fd_sc_hd__nor4_1 _11886_ (.A(_04557_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .D(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .Y(_05015_));
 sky130_fd_sc_hd__nor2_1 _11887_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__xnor2_1 _11888_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__nor2_1 _11889_ (.A(_05014_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__and2_1 _11890_ (.A(_05014_),
    .B(_05017_),
    .X(_05019_));
 sky130_fd_sc_hd__or2_1 _11891_ (.A(_05018_),
    .B(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__nor2_1 _11892_ (.A(_05013_),
    .B(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _11893_ (.A(_05013_),
    .B(_05020_),
    .Y(_05022_));
 sky130_fd_sc_hd__and2b_1 _11894_ (.A_N(_05021_),
    .B(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__or2_1 _11895_ (.A(_04765_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_05024_));
 sky130_fd_sc_hd__o211a_1 _11896_ (.A1(_04862_),
    .A2(_05023_),
    .B1(_05024_),
    .C1(_04739_),
    .X(_00635_));
 sky130_fd_sc_hd__or4_1 _11897_ (.A(_04557_),
    .B(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .C(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .D(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_05025_));
 sky130_fd_sc_hd__o21a_1 _11898_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_05025_),
    .B1(_04795_),
    .X(_05026_));
 sky130_fd_sc_hd__xor2_1 _11899_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__nand2_1 _11900_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__or2_1 _11901_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_05027_),
    .X(_05029_));
 sky130_fd_sc_hd__nand2_1 _11902_ (.A(_05028_),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__o21a_1 _11903_ (.A1(_05018_),
    .A2(_05021_),
    .B1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__o31ai_1 _11904_ (.A1(_05018_),
    .A2(_05021_),
    .A3(_05030_),
    .B1(_04758_),
    .Y(_05032_));
 sky130_fd_sc_hd__o221a_1 _11905_ (.A1(_04771_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B1(_05031_),
    .B2(_05032_),
    .C1(_04965_),
    .X(_00636_));
 sky130_fd_sc_hd__inv_2 _11906_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_05033_));
 sky130_fd_sc_hd__a21oi_1 _11907_ (.A1(_04952_),
    .A2(net114),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_05034_));
 sky130_fd_sc_hd__xnor2_1 _11908_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__or2_1 _11909_ (.A(_05033_),
    .B(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__nand2_1 _11910_ (.A(_05033_),
    .B(_05035_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _11911_ (.A(_05036_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__o21ai_1 _11912_ (.A1(_05014_),
    .A2(_05017_),
    .B1(_05028_),
    .Y(_05039_));
 sky130_fd_sc_hd__o21a_1 _11913_ (.A1(_05021_),
    .A2(_05039_),
    .B1(_05029_),
    .X(_05040_));
 sky130_fd_sc_hd__xnor2_1 _11914_ (.A(_05038_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_05041_),
    .S(_04757_),
    .X(_05042_));
 sky130_fd_sc_hd__and2_1 _11916_ (.A(_04850_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _11917_ (.A(_05043_),
    .X(_00637_));
 sky130_fd_sc_hd__inv_2 _11918_ (.A(_05038_),
    .Y(_05044_));
 sky130_fd_sc_hd__nand2_1 _11919_ (.A(_05044_),
    .B(_05040_),
    .Y(_05045_));
 sky130_fd_sc_hd__inv_2 _11920_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .Y(_05046_));
 sky130_fd_sc_hd__a31o_1 _11921_ (.A1(_05046_),
    .A2(_04952_),
    .A3(net114),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05047_));
 sky130_fd_sc_hd__xnor2_1 _11922_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__nand2_1 _11923_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__nor2_1 _11924_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_05048_),
    .Y(_05050_));
 sky130_fd_sc_hd__inv_2 _11925_ (.A(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__and2_1 _11926_ (.A(_05049_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__a21oi_1 _11927_ (.A1(_05036_),
    .A2(_05045_),
    .B1(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__a31o_1 _11928_ (.A1(_05036_),
    .A2(_05045_),
    .A3(_05052_),
    .B1(_04755_),
    .X(_05054_));
 sky130_fd_sc_hd__o221a_1 _11929_ (.A1(_04771_),
    .A2(net533),
    .B1(_05053_),
    .B2(_05054_),
    .C1(_04965_),
    .X(_00638_));
 sky130_fd_sc_hd__a21oi_1 _11930_ (.A1(_05036_),
    .A2(_05049_),
    .B1(_05050_),
    .Y(_05055_));
 sky130_fd_sc_hd__a41oi_2 _11931_ (.A1(_05029_),
    .A2(_05044_),
    .A3(_05039_),
    .A4(_05052_),
    .B1(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__nor2_1 _11932_ (.A(_05020_),
    .B(_05030_),
    .Y(_05057_));
 sky130_fd_sc_hd__o2111ai_2 _11933_ (.A1(_05005_),
    .A2(_05009_),
    .B1(_05044_),
    .C1(_05057_),
    .D1(_05052_),
    .Y(_05058_));
 sky130_fd_sc_hd__or2_1 _11934_ (.A(_04970_),
    .B(_05025_),
    .X(_05059_));
 sky130_fd_sc_hd__and2_1 _11935_ (.A(_04795_),
    .B(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__xnor2_1 _11936_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__nor2_1 _11937_ (.A(_04831_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__and2_1 _11938_ (.A(_04831_),
    .B(_05061_),
    .X(_05063_));
 sky130_fd_sc_hd__or2_1 _11939_ (.A(_05062_),
    .B(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__a21oi_1 _11940_ (.A1(_05056_),
    .A2(_05058_),
    .B1(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__and3_1 _11941_ (.A(_05064_),
    .B(_05056_),
    .C(_05058_),
    .X(_05066_));
 sky130_fd_sc_hd__nor2_1 _11942_ (.A(_05065_),
    .B(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__or2_1 _11943_ (.A(_04770_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_05068_));
 sky130_fd_sc_hd__o211a_1 _11944_ (.A1(_04862_),
    .A2(_05067_),
    .B1(_05068_),
    .C1(_04739_),
    .X(_00639_));
 sky130_fd_sc_hd__nor2_1 _11945_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05059_),
    .Y(_05069_));
 sky130_fd_sc_hd__nor2_1 _11946_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(_05070_),
    .A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .S(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_05071_));
 sky130_fd_sc_hd__buf_2 _11948_ (.A(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__and2_1 _11949_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_05069_),
    .X(_05073_));
 sky130_fd_sc_hd__o21a_1 _11950_ (.A1(_05072_),
    .A2(_05073_),
    .B1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_05074_));
 sky130_fd_sc_hd__or3_1 _11951_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_05072_),
    .C(_05073_),
    .X(_05075_));
 sky130_fd_sc_hd__and2b_1 _11952_ (.A_N(_05074_),
    .B(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(_05062_),
    .B(_05065_),
    .Y(_05077_));
 sky130_fd_sc_hd__xnor2_1 _11954_ (.A(_05076_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__or2_1 _11955_ (.A(_04770_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_4 _11956_ (.A(_04455_),
    .X(_05080_));
 sky130_fd_sc_hd__o211a_1 _11957_ (.A1(_04862_),
    .A2(_05078_),
    .B1(_05079_),
    .C1(_05080_),
    .X(_00640_));
 sky130_fd_sc_hd__clkbuf_4 _11958_ (.A(_05072_),
    .X(_05081_));
 sky130_fd_sc_hd__xor2_1 _11959_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__o31a_1 _11960_ (.A1(_05062_),
    .A2(_05065_),
    .A3(_05074_),
    .B1(_05075_),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_1 _11961_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__and2_1 _11962_ (.A(_05082_),
    .B(_05083_),
    .X(_05085_));
 sky130_fd_sc_hd__o21ai_1 _11963_ (.A1(_05084_),
    .A2(_05085_),
    .B1(_04786_),
    .Y(_05086_));
 sky130_fd_sc_hd__o211a_1 _11964_ (.A1(_04769_),
    .A2(net545),
    .B1(_04979_),
    .C1(_05086_),
    .X(_00641_));
 sky130_fd_sc_hd__xor2_1 _11965_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_05081_),
    .X(_05087_));
 sky130_fd_sc_hd__a21oi_1 _11966_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(_05081_),
    .B1(_05085_),
    .Y(_05088_));
 sky130_fd_sc_hd__and2_1 _11967_ (.A(_05087_),
    .B(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__o21ai_1 _11968_ (.A1(_05087_),
    .A2(_05088_),
    .B1(_04786_),
    .Y(_05090_));
 sky130_fd_sc_hd__o221a_1 _11969_ (.A1(_04771_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_05089_),
    .B2(_05090_),
    .C1(_04965_),
    .X(_00642_));
 sky130_fd_sc_hd__o21a_1 _11970_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_05081_),
    .X(_05091_));
 sky130_fd_sc_hd__a31o_1 _11971_ (.A1(_05082_),
    .A2(_05083_),
    .A3(_05087_),
    .B1(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__or2_1 _11972_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05072_),
    .X(_05093_));
 sky130_fd_sc_hd__nand2_1 _11973_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05072_),
    .Y(_05094_));
 sky130_fd_sc_hd__and2_1 _11974_ (.A(_05093_),
    .B(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__xor2_1 _11975_ (.A(_05092_),
    .B(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__or2_1 _11976_ (.A(_04770_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_05097_));
 sky130_fd_sc_hd__o211a_1 _11977_ (.A1(_04862_),
    .A2(_05096_),
    .B1(_05097_),
    .C1(_05080_),
    .X(_00643_));
 sky130_fd_sc_hd__a21bo_1 _11978_ (.A1(_05092_),
    .A2(_05095_),
    .B1_N(_05094_),
    .X(_05098_));
 sky130_fd_sc_hd__xor2_1 _11979_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_05072_),
    .X(_05099_));
 sky130_fd_sc_hd__xor2_1 _11980_ (.A(_05098_),
    .B(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__or2_1 _11981_ (.A(_04770_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_05101_));
 sky130_fd_sc_hd__o211a_1 _11982_ (.A1(_04862_),
    .A2(_05100_),
    .B1(_05101_),
    .C1(_05080_),
    .X(_00644_));
 sky130_fd_sc_hd__nor2_1 _11983_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05072_),
    .Y(_05102_));
 sky130_fd_sc_hd__and2_1 _11984_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05072_),
    .X(_05103_));
 sky130_fd_sc_hd__nor2_1 _11985_ (.A(_05102_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__and2_1 _11986_ (.A(_05095_),
    .B(_05099_),
    .X(_05105_));
 sky130_fd_sc_hd__o21a_1 _11987_ (.A1(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_05081_),
    .X(_05106_));
 sky130_fd_sc_hd__a21oi_1 _11988_ (.A1(_05092_),
    .A2(_05105_),
    .B1(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__xnor2_1 _11989_ (.A(_05104_),
    .B(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__mux2_1 _11990_ (.A0(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A1(_05108_),
    .S(_04757_),
    .X(_05109_));
 sky130_fd_sc_hd__and2_1 _11991_ (.A(_04850_),
    .B(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__clkbuf_1 _11992_ (.A(_05110_),
    .X(_00645_));
 sky130_fd_sc_hd__o21ba_1 _11993_ (.A1(_05102_),
    .A2(_05107_),
    .B1_N(_05103_),
    .X(_05111_));
 sky130_fd_sc_hd__xor2_1 _11994_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_05081_),
    .X(_05112_));
 sky130_fd_sc_hd__and2_1 _11995_ (.A(_05111_),
    .B(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__o21ai_1 _11996_ (.A1(_05111_),
    .A2(_05112_),
    .B1(_04786_),
    .Y(_05114_));
 sky130_fd_sc_hd__o221a_1 _11997_ (.A1(_04771_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_05113_),
    .B2(_05114_),
    .C1(_04965_),
    .X(_00646_));
 sky130_fd_sc_hd__or2_1 _11998_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05081_),
    .X(_05115_));
 sky130_fd_sc_hd__nand2_1 _11999_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05081_),
    .Y(_05116_));
 sky130_fd_sc_hd__and2_1 _12000_ (.A(_05115_),
    .B(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__and3_1 _12001_ (.A(_05104_),
    .B(_05105_),
    .C(_05112_),
    .X(_05118_));
 sky130_fd_sc_hd__a22o_1 _12002_ (.A1(_04903_),
    .A2(_05081_),
    .B1(_05092_),
    .B2(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__nand2_1 _12003_ (.A(_05117_),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__o21a_1 _12004_ (.A1(_05117_),
    .A2(_05119_),
    .B1(_04757_),
    .X(_05121_));
 sky130_fd_sc_hd__a22o_1 _12005_ (.A1(_04754_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B1(_05120_),
    .B2(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__and2_1 _12006_ (.A(_04850_),
    .B(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_1 _12007_ (.A(_05123_),
    .X(_00647_));
 sky130_fd_sc_hd__xor2_1 _12008_ (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05081_),
    .X(_05124_));
 sky130_fd_sc_hd__a21oi_1 _12009_ (.A1(_05116_),
    .A2(_05120_),
    .B1(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__a31o_1 _12010_ (.A1(_05116_),
    .A2(_05120_),
    .A3(_05124_),
    .B1(_04754_),
    .X(_05126_));
 sky130_fd_sc_hd__o221a_1 _12011_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_04769_),
    .B1(_05125_),
    .B2(_05126_),
    .C1(_04965_),
    .X(_00648_));
 sky130_fd_sc_hd__and2_1 _12012_ (.A(_04758_),
    .B(_02310_),
    .X(_05127_));
 sky130_fd_sc_hd__clkbuf_1 _12013_ (.A(_05127_),
    .X(_00649_));
 sky130_fd_sc_hd__inv_2 _12014_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_05128_));
 sky130_fd_sc_hd__clkbuf_4 _12015_ (.A(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__clkbuf_4 _12016_ (.A(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__or2_1 _12017_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_01250_),
    .X(_05131_));
 sky130_fd_sc_hd__o211a_1 _12018_ (.A1(_05130_),
    .A2(net183),
    .B1(_04979_),
    .C1(_05131_),
    .X(_00650_));
 sky130_fd_sc_hd__clkbuf_4 _12019_ (.A(_01249_),
    .X(_05132_));
 sky130_fd_sc_hd__or2_1 _12020_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__o211a_1 _12021_ (.A1(_05130_),
    .A2(net218),
    .B1(_04979_),
    .C1(_05133_),
    .X(_00651_));
 sky130_fd_sc_hd__or2_1 _12022_ (.A(net149),
    .B(_05132_),
    .X(_05134_));
 sky130_fd_sc_hd__o211a_1 _12023_ (.A1(_05130_),
    .A2(net257),
    .B1(_04979_),
    .C1(_05134_),
    .X(_00652_));
 sky130_fd_sc_hd__or2_1 _12024_ (.A(net153),
    .B(_05132_),
    .X(_05135_));
 sky130_fd_sc_hd__o211a_1 _12025_ (.A1(_05130_),
    .A2(net209),
    .B1(_04979_),
    .C1(_05135_),
    .X(_00653_));
 sky130_fd_sc_hd__or2_1 _12026_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(_05132_),
    .X(_05136_));
 sky130_fd_sc_hd__o211a_1 _12027_ (.A1(_05130_),
    .A2(net162),
    .B1(_04979_),
    .C1(_05136_),
    .X(_00654_));
 sky130_fd_sc_hd__or2_1 _12028_ (.A(net169),
    .B(_05132_),
    .X(_05137_));
 sky130_fd_sc_hd__o211a_1 _12029_ (.A1(_05130_),
    .A2(net205),
    .B1(_04979_),
    .C1(_05137_),
    .X(_00655_));
 sky130_fd_sc_hd__or2_1 _12030_ (.A(_01250_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(_05138_));
 sky130_fd_sc_hd__o211a_1 _12031_ (.A1(_05130_),
    .A2(net201),
    .B1(_04979_),
    .C1(_05138_),
    .X(_00656_));
 sky130_fd_sc_hd__buf_2 _12032_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05139_));
 sky130_fd_sc_hd__buf_4 _12033_ (.A(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__buf_4 _12034_ (.A(_03619_),
    .X(_05141_));
 sky130_fd_sc_hd__buf_4 _12035_ (.A(_05139_),
    .X(_05142_));
 sky130_fd_sc_hd__nand2_1 _12036_ (.A(_05142_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .Y(_05143_));
 sky130_fd_sc_hd__o211a_1 _12037_ (.A1(_05140_),
    .A2(net342),
    .B1(_05141_),
    .C1(_05143_),
    .X(_00657_));
 sky130_fd_sc_hd__nand2_1 _12038_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .Y(_05144_));
 sky130_fd_sc_hd__or2_1 _12039_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(_05145_));
 sky130_fd_sc_hd__a21oi_1 _12040_ (.A1(_05144_),
    .A2(_05145_),
    .B1(_04829_),
    .Y(_05146_));
 sky130_fd_sc_hd__a31o_1 _12041_ (.A1(_04829_),
    .A2(_05144_),
    .A3(_05145_),
    .B1(_05129_),
    .X(_05147_));
 sky130_fd_sc_hd__o221a_1 _12042_ (.A1(_05140_),
    .A2(net507),
    .B1(_05146_),
    .B2(_05147_),
    .C1(_04965_),
    .X(_00658_));
 sky130_fd_sc_hd__and3_1 _12043_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(_05148_));
 sky130_fd_sc_hd__a21oi_1 _12044_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_05149_));
 sky130_fd_sc_hd__or2_1 _12045_ (.A(_05148_),
    .B(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__nor2_1 _12046_ (.A(_05146_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__a21o_1 _12047_ (.A1(_05146_),
    .A2(_05150_),
    .B1(_05129_),
    .X(_05152_));
 sky130_fd_sc_hd__o221a_1 _12048_ (.A1(_05140_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B1(_05151_),
    .B2(_05152_),
    .C1(_04965_),
    .X(_00659_));
 sky130_fd_sc_hd__clkbuf_4 _12049_ (.A(_05139_),
    .X(_05153_));
 sky130_fd_sc_hd__nand2_1 _12050_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05148_),
    .Y(_05154_));
 sky130_fd_sc_hd__o31a_1 _12051_ (.A1(_04829_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A3(_05145_),
    .B1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__and2_1 _12052_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__o21ai_1 _12053_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_05155_),
    .B1(_01250_),
    .Y(_05157_));
 sky130_fd_sc_hd__o221a_1 _12054_ (.A1(_05153_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B1(_05156_),
    .B2(_05157_),
    .C1(_04965_),
    .X(_00660_));
 sky130_fd_sc_hd__or3_1 _12055_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .C(_05145_),
    .X(_05158_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_05148_),
    .Y(_05159_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(_05158_),
    .A1(_05159_),
    .S(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05160_));
 sky130_fd_sc_hd__and2_1 _12058_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__o21ai_1 _12059_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_05160_),
    .B1(_01250_),
    .Y(_05162_));
 sky130_fd_sc_hd__o221a_1 _12060_ (.A1(_05153_),
    .A2(net525),
    .B1(_05161_),
    .B2(_05162_),
    .C1(_04965_),
    .X(_00661_));
 sky130_fd_sc_hd__inv_2 _12061_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_05163_));
 sky130_fd_sc_hd__clkbuf_4 _12062_ (.A(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__o21ai_1 _12063_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_05158_),
    .B1(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__a31o_1 _12064_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A3(_05148_),
    .B1(_05164_),
    .X(_05166_));
 sky130_fd_sc_hd__inv_2 _12065_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .Y(_05167_));
 sky130_fd_sc_hd__a21oi_1 _12066_ (.A1(_05165_),
    .A2(_05166_),
    .B1(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__a31o_1 _12067_ (.A1(_05167_),
    .A2(_05165_),
    .A3(_05166_),
    .B1(_05129_),
    .X(_05169_));
 sky130_fd_sc_hd__clkbuf_4 _12068_ (.A(_04538_),
    .X(_05170_));
 sky130_fd_sc_hd__o221a_1 _12069_ (.A1(_05153_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_05168_),
    .B2(_05169_),
    .C1(_05170_),
    .X(_00662_));
 sky130_fd_sc_hd__and4_1 _12070_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .D(_05148_),
    .X(_05171_));
 sky130_fd_sc_hd__or3_1 _12071_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(_05158_),
    .X(_05172_));
 sky130_fd_sc_hd__inv_2 _12072_ (.A(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__mux2_1 _12073_ (.A0(_05171_),
    .A1(_05173_),
    .S(_05164_),
    .X(_05174_));
 sky130_fd_sc_hd__xnor2_1 _12074_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_1 _12075_ (.A(_05142_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__o211a_1 _12076_ (.A1(_05140_),
    .A2(net643),
    .B1(_05141_),
    .C1(_05176_),
    .X(_00663_));
 sky130_fd_sc_hd__or2_1 _12077_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_05172_),
    .X(_05177_));
 sky130_fd_sc_hd__nor2_1 _12078_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a31o_1 _12079_ (.A1(_04829_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(_05171_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__xor2_1 _12080_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__or2_1 _12081_ (.A(_05132_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(_05181_));
 sky130_fd_sc_hd__o211a_1 _12082_ (.A1(_05130_),
    .A2(_05180_),
    .B1(_05181_),
    .C1(_05080_),
    .X(_00664_));
 sky130_fd_sc_hd__and3_1 _12083_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_05171_),
    .X(_05182_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__o31a_1 _12085_ (.A1(_04829_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A3(_05177_),
    .B1(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__and2_1 _12086_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__o21ai_1 _12087_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_05184_),
    .B1(_01250_),
    .Y(_05186_));
 sky130_fd_sc_hd__o221a_1 _12088_ (.A1(_05153_),
    .A2(net529),
    .B1(_05185_),
    .B2(_05186_),
    .C1(_05170_),
    .X(_00665_));
 sky130_fd_sc_hd__nand3_1 _12089_ (.A(_04829_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_05182_),
    .Y(_05187_));
 sky130_fd_sc_hd__o41a_1 _12090_ (.A1(_04829_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A3(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A4(_05177_),
    .B1(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__nor2_1 _12091_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__a21o_1 _12092_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_05188_),
    .B1(_05129_),
    .X(_05190_));
 sky130_fd_sc_hd__o221a_1 _12093_ (.A1(_05153_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_05189_),
    .B2(_05190_),
    .C1(_05170_),
    .X(_00666_));
 sky130_fd_sc_hd__or4_1 _12094_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .D(_05177_),
    .X(_05191_));
 sky130_fd_sc_hd__and3_1 _12095_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_05182_),
    .X(_05192_));
 sky130_fd_sc_hd__nand2_1 _12096_ (.A(_04829_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__o21a_1 _12097_ (.A1(_04829_),
    .A2(_05191_),
    .B1(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__and2_1 _12098_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__o21ai_1 _12099_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05194_),
    .B1(_01250_),
    .Y(_05196_));
 sky130_fd_sc_hd__o221a_1 _12100_ (.A1(_05153_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_05195_),
    .B2(_05196_),
    .C1(_05170_),
    .X(_00667_));
 sky130_fd_sc_hd__o21a_1 _12101_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05191_),
    .B1(_05164_),
    .X(_05197_));
 sky130_fd_sc_hd__a21o_1 _12102_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05192_),
    .B1(_05164_),
    .X(_05198_));
 sky130_fd_sc_hd__or2b_1 _12103_ (.A(_05197_),
    .B_N(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__nor2_1 _12104_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__a21o_1 _12105_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_05199_),
    .B1(_05129_),
    .X(_05201_));
 sky130_fd_sc_hd__o221a_1 _12106_ (.A1(_05153_),
    .A2(net485),
    .B1(_05200_),
    .B2(_05201_),
    .C1(_05170_),
    .X(_00668_));
 sky130_fd_sc_hd__a21oi_1 _12107_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_05198_),
    .B1(_05197_),
    .Y(_05202_));
 sky130_fd_sc_hd__buf_2 _12108_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05203_));
 sky130_fd_sc_hd__or2_1 _12109_ (.A(_05132_),
    .B(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__o211a_1 _12110_ (.A1(_05130_),
    .A2(_05202_),
    .B1(_05204_),
    .C1(_05080_),
    .X(_00669_));
 sky130_fd_sc_hd__inv_2 _12111_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .Y(_05205_));
 sky130_fd_sc_hd__nor2_1 _12112_ (.A(_05205_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_05206_));
 sky130_fd_sc_hd__a21o_1 _12113_ (.A1(_05205_),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_05129_),
    .X(_05207_));
 sky130_fd_sc_hd__o221a_1 _12114_ (.A1(_05153_),
    .A2(net424),
    .B1(_05206_),
    .B2(_05207_),
    .C1(_05170_),
    .X(_00670_));
 sky130_fd_sc_hd__and2b_1 _12115_ (.A_N(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_05208_));
 sky130_fd_sc_hd__xnor2_1 _12116_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__xnor2_1 _12117_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__xor2_1 _12118_ (.A(_05206_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__or2_1 _12119_ (.A(_05132_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_05212_));
 sky130_fd_sc_hd__o211a_1 _12120_ (.A1(_05130_),
    .A2(_05211_),
    .B1(_05212_),
    .C1(_05080_),
    .X(_00671_));
 sky130_fd_sc_hd__o21a_1 _12121_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_05163_),
    .X(_05213_));
 sky130_fd_sc_hd__xnor2_1 _12122_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__nor2_1 _12123_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_1 _12124_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_05214_),
    .Y(_05216_));
 sky130_fd_sc_hd__or2b_1 _12125_ (.A(_05215_),
    .B_N(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__nand2_1 _12126_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_05209_),
    .Y(_05218_));
 sky130_fd_sc_hd__o21a_1 _12127_ (.A1(_05206_),
    .A2(_05210_),
    .B1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__a21o_1 _12128_ (.A1(_05217_),
    .A2(_05219_),
    .B1(_05128_),
    .X(_05220_));
 sky130_fd_sc_hd__nor2_1 _12129_ (.A(_05217_),
    .B(_05219_),
    .Y(_05221_));
 sky130_fd_sc_hd__clkbuf_4 _12130_ (.A(_05128_),
    .X(_05222_));
 sky130_fd_sc_hd__a2bb2o_1 _12131_ (.A1_N(_05220_),
    .A2_N(_05221_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B2(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__and2_1 _12132_ (.A(_04850_),
    .B(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__clkbuf_1 _12133_ (.A(_05224_),
    .X(_00672_));
 sky130_fd_sc_hd__o31a_1 _12134_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_05163_),
    .X(_05225_));
 sky130_fd_sc_hd__xnor2_1 _12135_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__and2_1 _12136_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__or2_1 _12137_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_05226_),
    .X(_05228_));
 sky130_fd_sc_hd__and2b_1 _12138_ (.A_N(_05227_),
    .B(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__o21ai_1 _12139_ (.A1(_05215_),
    .A2(_05219_),
    .B1(_05216_),
    .Y(_05230_));
 sky130_fd_sc_hd__xor2_1 _12140_ (.A(_05229_),
    .B(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_05231_),
    .S(_01249_),
    .X(_05232_));
 sky130_fd_sc_hd__and2_1 _12142_ (.A(_04850_),
    .B(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _12143_ (.A(_05233_),
    .X(_00673_));
 sky130_fd_sc_hd__clkbuf_4 _12144_ (.A(_05222_),
    .X(_05234_));
 sky130_fd_sc_hd__a21o_1 _12145_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_05227_),
    .X(_05235_));
 sky130_fd_sc_hd__or4_4 _12146_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .D(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_05236_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_05163_),
    .B(net121),
    .Y(_05237_));
 sky130_fd_sc_hd__xor2_1 _12148_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__and2_1 _12149_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__nor2_1 _12150_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_05238_),
    .Y(_05240_));
 sky130_fd_sc_hd__nor2_1 _12151_ (.A(_05239_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__xor2_1 _12152_ (.A(_05235_),
    .B(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__or2_1 _12153_ (.A(_05132_),
    .B(net482),
    .X(_05243_));
 sky130_fd_sc_hd__o211a_1 _12154_ (.A1(_05234_),
    .A2(_05242_),
    .B1(_05243_),
    .C1(_05080_),
    .X(_00674_));
 sky130_fd_sc_hd__o21a_1 _12155_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(net121),
    .B1(_05163_),
    .X(_05244_));
 sky130_fd_sc_hd__xor2_1 _12156_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__nand2b_2 _12157_ (.A_N(_05245_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .Y(_05246_));
 sky130_fd_sc_hd__or2b_1 _12158_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B_N(_05245_),
    .X(_05247_));
 sky130_fd_sc_hd__nand2_1 _12159_ (.A(_05246_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__a21o_1 _12160_ (.A1(_05235_),
    .A2(_05241_),
    .B1(_05239_),
    .X(_05249_));
 sky130_fd_sc_hd__and2_1 _12161_ (.A(_05248_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__o21ai_1 _12162_ (.A1(_05248_),
    .A2(_05249_),
    .B1(_01250_),
    .Y(_05251_));
 sky130_fd_sc_hd__o221a_1 _12163_ (.A1(_05153_),
    .A2(net484),
    .B1(_05250_),
    .B2(_05251_),
    .C1(_05170_),
    .X(_00675_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(_05247_),
    .B(_05249_),
    .Y(_05252_));
 sky130_fd_sc_hd__o31a_1 _12165_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A3(net121),
    .B1(_05163_),
    .X(_05253_));
 sky130_fd_sc_hd__xnor2_2 _12166_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__xnor2_2 _12167_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__a21o_1 _12168_ (.A1(_05246_),
    .A2(_05252_),
    .B1(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__a31oi_1 _12169_ (.A1(_05246_),
    .A2(_05252_),
    .A3(_05255_),
    .B1(_05128_),
    .Y(_05257_));
 sky130_fd_sc_hd__a22o_1 _12170_ (.A1(_05222_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_05256_),
    .B2(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__and2_1 _12171_ (.A(_04850_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__clkbuf_1 _12172_ (.A(_05259_),
    .X(_00676_));
 sky130_fd_sc_hd__or4_4 _12173_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .D(_05236_),
    .X(_05260_));
 sky130_fd_sc_hd__and2_4 _12174_ (.A(_05260_),
    .B(_05163_),
    .X(_05261_));
 sky130_fd_sc_hd__xnor2_1 _12175_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__and2_4 _12176_ (.A(_05262_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_05263_));
 sky130_fd_sc_hd__nor2_1 _12177_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_05262_),
    .Y(_05264_));
 sky130_fd_sc_hd__or2_4 _12178_ (.A(_05263_),
    .B(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__a21bo_1 _12179_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(_05254_),
    .B1_N(_05256_),
    .X(_05266_));
 sky130_fd_sc_hd__xnor2_1 _12180_ (.A(_05265_),
    .B(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__or2_1 _12181_ (.A(_05132_),
    .B(net517),
    .X(_05268_));
 sky130_fd_sc_hd__o211a_1 _12182_ (.A1(_05234_),
    .A2(_05267_),
    .B1(_05268_),
    .C1(_05080_),
    .X(_00677_));
 sky130_fd_sc_hd__inv_2 _12183_ (.A(_05246_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_1 _12184_ (.A1(_05239_),
    .A2(_05269_),
    .B1(_05247_),
    .Y(_05270_));
 sky130_fd_sc_hd__a21oi_1 _12185_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(_05254_),
    .B1(_05263_),
    .Y(_05271_));
 sky130_fd_sc_hd__o32a_1 _12186_ (.A1(_05255_),
    .A2(_05270_),
    .A3(_05265_),
    .B1(_05271_),
    .B2(_05264_),
    .X(_05272_));
 sky130_fd_sc_hd__nand3_1 _12187_ (.A(_05241_),
    .B(_05246_),
    .C(_05247_),
    .Y(_05273_));
 sky130_fd_sc_hd__or4b_4 _12188_ (.A(_05255_),
    .B(_05273_),
    .C(_05265_),
    .D_N(_05235_),
    .X(_05274_));
 sky130_fd_sc_hd__inv_2 _12189_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_05275_));
 sky130_fd_sc_hd__or2_1 _12190_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05260_),
    .X(_05276_));
 sky130_fd_sc_hd__a21oi_1 _12191_ (.A1(_05163_),
    .A2(_05276_),
    .B1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_05277_));
 sky130_fd_sc_hd__a21o_1 _12192_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_05164_),
    .B1(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_4 _12193_ (.A(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__o21a_1 _12194_ (.A1(_05275_),
    .A2(_05276_),
    .B1(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__xnor2_1 _12195_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__a21o_1 _12196_ (.A1(_05272_),
    .A2(_05274_),
    .B1(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__nand3_1 _12197_ (.A(_05281_),
    .B(_05272_),
    .C(_05274_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21o_1 _12198_ (.A1(_05282_),
    .A2(_05283_),
    .B1(_05234_),
    .X(_05284_));
 sky130_fd_sc_hd__o211a_1 _12199_ (.A1(_05140_),
    .A2(net640),
    .B1(_05141_),
    .C1(_05284_),
    .X(_00678_));
 sky130_fd_sc_hd__xnor2_1 _12200_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_05279_),
    .Y(_05285_));
 sky130_fd_sc_hd__and2_1 _12201_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_05280_),
    .X(_05286_));
 sky130_fd_sc_hd__or2b_1 _12202_ (.A(_05286_),
    .B_N(_05282_),
    .X(_05287_));
 sky130_fd_sc_hd__xnor2_1 _12203_ (.A(_05285_),
    .B(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__or2_1 _12204_ (.A(_05139_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_05289_));
 sky130_fd_sc_hd__o211a_1 _12205_ (.A1(_05234_),
    .A2(_05288_),
    .B1(_05289_),
    .C1(_05080_),
    .X(_00679_));
 sky130_fd_sc_hd__buf_2 _12206_ (.A(_01252_),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_4 _12207_ (.A(_05279_),
    .X(_05291_));
 sky130_fd_sc_hd__a21o_1 _12208_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_05291_),
    .B1(_05286_),
    .X(_05292_));
 sky130_fd_sc_hd__o21ba_1 _12209_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_05291_),
    .B1_N(_05282_),
    .X(_05293_));
 sky130_fd_sc_hd__nor2_1 _12210_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_05279_),
    .Y(_05294_));
 sky130_fd_sc_hd__and2_1 _12211_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_05279_),
    .X(_05295_));
 sky130_fd_sc_hd__or2_1 _12212_ (.A(_05294_),
    .B(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__or3b_1 _12213_ (.A(_05292_),
    .B(_05293_),
    .C_N(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_01249_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21ba_1 _12215_ (.A1(_05292_),
    .A2(_05293_),
    .B1_N(_05296_),
    .X(_05299_));
 sky130_fd_sc_hd__a2bb2o_1 _12216_ (.A1_N(_05298_),
    .A2_N(_05299_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B2(_05128_),
    .X(_05300_));
 sky130_fd_sc_hd__and2_1 _12217_ (.A(_05290_),
    .B(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__clkbuf_1 _12218_ (.A(_05301_),
    .X(_00680_));
 sky130_fd_sc_hd__xnor2_1 _12219_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_05279_),
    .Y(_05302_));
 sky130_fd_sc_hd__o21a_1 _12220_ (.A1(_05295_),
    .A2(_05299_),
    .B1(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__o31ai_1 _12221_ (.A1(_05295_),
    .A2(_05299_),
    .A3(_05302_),
    .B1(_01250_),
    .Y(_05304_));
 sky130_fd_sc_hd__o221a_1 _12222_ (.A1(_05153_),
    .A2(net570),
    .B1(_05303_),
    .B2(_05304_),
    .C1(_05170_),
    .X(_00681_));
 sky130_fd_sc_hd__or2_1 _12223_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05279_),
    .X(_05305_));
 sky130_fd_sc_hd__nand2_1 _12224_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05279_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_1 _12225_ (.A(_05305_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__or4_4 _12226_ (.A(_05282_),
    .B(_05285_),
    .C(_05296_),
    .D(_05302_),
    .X(_05308_));
 sky130_fd_sc_hd__a211oi_1 _12227_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(_05291_),
    .B1(_05295_),
    .C1(_05292_),
    .Y(_05309_));
 sky130_fd_sc_hd__and2_1 _12228_ (.A(_05308_),
    .B(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__xor2_1 _12229_ (.A(_05307_),
    .B(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__or2_1 _12230_ (.A(_05139_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_05312_));
 sky130_fd_sc_hd__o211a_1 _12231_ (.A1(_05234_),
    .A2(_05311_),
    .B1(_05312_),
    .C1(_05080_),
    .X(_00682_));
 sky130_fd_sc_hd__xnor2_1 _12232_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_05279_),
    .Y(_05313_));
 sky130_fd_sc_hd__o21ai_1 _12233_ (.A1(_05307_),
    .A2(_05310_),
    .B1(_05306_),
    .Y(_05314_));
 sky130_fd_sc_hd__nor2_1 _12234_ (.A(_05313_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__a21o_1 _12235_ (.A1(_05313_),
    .A2(_05314_),
    .B1(_05129_),
    .X(_05316_));
 sky130_fd_sc_hd__o221a_1 _12236_ (.A1(_05142_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_05315_),
    .B2(_05316_),
    .C1(_05170_),
    .X(_00683_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_05279_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _12238_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_05291_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _12239_ (.A(_05317_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__or2_1 _12240_ (.A(_05307_),
    .B(_05313_),
    .X(_05320_));
 sky130_fd_sc_hd__o21ai_1 _12241_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_05291_),
    .Y(_05321_));
 sky130_fd_sc_hd__o21a_1 _12242_ (.A1(_05310_),
    .A2(_05320_),
    .B1(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__xor2_1 _12243_ (.A(_05319_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A1(_05323_),
    .S(_01249_),
    .X(_05324_));
 sky130_fd_sc_hd__and2_1 _12245_ (.A(_05290_),
    .B(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _12246_ (.A(_05325_),
    .X(_00684_));
 sky130_fd_sc_hd__xnor2_1 _12247_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_05291_),
    .Y(_05326_));
 sky130_fd_sc_hd__o21ai_1 _12248_ (.A1(_05319_),
    .A2(_05322_),
    .B1(_05318_),
    .Y(_05327_));
 sky130_fd_sc_hd__nor2_1 _12249_ (.A(_05326_),
    .B(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__a21o_1 _12250_ (.A1(_05326_),
    .A2(_05327_),
    .B1(_05129_),
    .X(_05329_));
 sky130_fd_sc_hd__o221a_1 _12251_ (.A1(_05142_),
    .A2(net594),
    .B1(_05328_),
    .B2(_05329_),
    .C1(_05170_),
    .X(_00685_));
 sky130_fd_sc_hd__or2_1 _12252_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05291_),
    .X(_05330_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05291_),
    .Y(_05331_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_05330_),
    .B(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__or4_4 _12255_ (.A(_05308_),
    .B(_05319_),
    .C(_05320_),
    .D(_05326_),
    .X(_05333_));
 sky130_fd_sc_hd__o21ai_1 _12256_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_05291_),
    .Y(_05334_));
 sky130_fd_sc_hd__and4_1 _12257_ (.A(_05309_),
    .B(_05321_),
    .C(_05333_),
    .D(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__xor2_1 _12258_ (.A(_05332_),
    .B(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A1(_05336_),
    .S(_01249_),
    .X(_05337_));
 sky130_fd_sc_hd__and2_1 _12260_ (.A(_05290_),
    .B(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_1 _12261_ (.A(_05338_),
    .X(_00686_));
 sky130_fd_sc_hd__o21ai_1 _12262_ (.A1(_05332_),
    .A2(_05335_),
    .B1(_05331_),
    .Y(_05339_));
 sky130_fd_sc_hd__xnor2_1 _12263_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_05291_),
    .Y(_05340_));
 sky130_fd_sc_hd__xnor2_1 _12264_ (.A(_05339_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__or2_1 _12265_ (.A(_05139_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_4 _12266_ (.A(_04455_),
    .X(_05343_));
 sky130_fd_sc_hd__o211a_1 _12267_ (.A1(_05234_),
    .A2(_05341_),
    .B1(_05342_),
    .C1(_05343_),
    .X(_00687_));
 sky130_fd_sc_hd__and2_1 _12268_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_05344_));
 sky130_fd_sc_hd__nor2_1 _12269_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .Y(_05345_));
 sky130_fd_sc_hd__o21ai_2 _12270_ (.A1(_05344_),
    .A2(_05345_),
    .B1(_05142_),
    .Y(_05346_));
 sky130_fd_sc_hd__o211a_1 _12271_ (.A1(_05140_),
    .A2(net272),
    .B1(_05141_),
    .C1(_05346_),
    .X(_00688_));
 sky130_fd_sc_hd__and2b_1 _12272_ (.A_N(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_05347_));
 sky130_fd_sc_hd__xnor2_1 _12273_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__xnor2_1 _12274_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nor2_1 _12275_ (.A(_05344_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__and2_1 _12276_ (.A(_05344_),
    .B(_05349_),
    .X(_05351_));
 sky130_fd_sc_hd__o21ai_2 _12277_ (.A1(_05350_),
    .A2(_05351_),
    .B1(_01250_),
    .Y(_05352_));
 sky130_fd_sc_hd__o211a_1 _12278_ (.A1(_05140_),
    .A2(net321),
    .B1(_05141_),
    .C1(_05352_),
    .X(_00689_));
 sky130_fd_sc_hd__and2b_1 _12279_ (.A_N(_05348_),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_05353_));
 sky130_fd_sc_hd__o21a_1 _12280_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_05164_),
    .X(_05354_));
 sky130_fd_sc_hd__xnor2_1 _12281_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__xnor2_1 _12282_ (.A(_04996_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__o21bai_2 _12283_ (.A1(_05353_),
    .A2(_05351_),
    .B1_N(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__or3b_1 _12284_ (.A(_05353_),
    .B(_05351_),
    .C_N(_05356_),
    .X(_05358_));
 sky130_fd_sc_hd__inv_2 _12285_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_05359_));
 sky130_fd_sc_hd__nor2_1 _12286_ (.A(_01249_),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__a31o_1 _12287_ (.A1(_05139_),
    .A2(_05357_),
    .A3(_05358_),
    .B1(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__and2_1 _12288_ (.A(_05290_),
    .B(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _12289_ (.A(_05362_),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _12290_ (.A(_04996_),
    .B(_05355_),
    .X(_05363_));
 sky130_fd_sc_hd__o31a_1 _12291_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A3(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_05164_),
    .X(_05364_));
 sky130_fd_sc_hd__xnor2_1 _12292_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__nor2_1 _12293_ (.A(_05000_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__and2_1 _12294_ (.A(_05000_),
    .B(_05365_),
    .X(_05367_));
 sky130_fd_sc_hd__or2_1 _12295_ (.A(_05366_),
    .B(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__and3_1 _12296_ (.A(_05363_),
    .B(_05357_),
    .C(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__a21oi_1 _12297_ (.A1(_05363_),
    .A2(_05357_),
    .B1(_05368_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_1 _12298_ (.A(_05128_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_05371_));
 sky130_fd_sc_hd__o31a_1 _12299_ (.A1(_05128_),
    .A2(_05369_),
    .A3(_05370_),
    .B1(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__and2b_1 _12300_ (.A_N(_05372_),
    .B(_03118_),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _12301_ (.A(_05373_),
    .X(_00691_));
 sky130_fd_sc_hd__or2_1 _12302_ (.A(_05366_),
    .B(_05370_),
    .X(_05374_));
 sky130_fd_sc_hd__or4_2 _12303_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .D(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_05375_));
 sky130_fd_sc_hd__nand2_1 _12304_ (.A(_05163_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__xor2_1 _12305_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__xnor2_1 _12306_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__nand2_1 _12307_ (.A(_05374_),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__or2_1 _12308_ (.A(_05374_),
    .B(_05378_),
    .X(_05380_));
 sky130_fd_sc_hd__a21o_1 _12309_ (.A1(_05379_),
    .A2(_05380_),
    .B1(_05234_),
    .X(_05381_));
 sky130_fd_sc_hd__o211a_1 _12310_ (.A1(_05140_),
    .A2(net289),
    .B1(_05141_),
    .C1(_05381_),
    .X(_00692_));
 sky130_fd_sc_hd__or2b_1 _12311_ (.A(_05377_),
    .B_N(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_05382_));
 sky130_fd_sc_hd__inv_2 _12312_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .Y(_05383_));
 sky130_fd_sc_hd__o21a_1 _12313_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(_05375_),
    .B1(_05164_),
    .X(_05384_));
 sky130_fd_sc_hd__xnor2_1 _12314_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__nor2_1 _12315_ (.A(_05383_),
    .B(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__and2_1 _12316_ (.A(_05383_),
    .B(_05385_),
    .X(_05387_));
 sky130_fd_sc_hd__nor2_1 _12317_ (.A(_05386_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__a21oi_1 _12318_ (.A1(_05382_),
    .A2(_05379_),
    .B1(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a31o_1 _12319_ (.A1(_05382_),
    .A2(_05379_),
    .A3(_05388_),
    .B1(_05222_),
    .X(_05390_));
 sky130_fd_sc_hd__clkbuf_4 _12320_ (.A(_04538_),
    .X(_05391_));
 sky130_fd_sc_hd__o221a_1 _12321_ (.A1(_05142_),
    .A2(net420),
    .B1(_05389_),
    .B2(_05390_),
    .C1(_05391_),
    .X(_00693_));
 sky130_fd_sc_hd__inv_2 _12322_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_05392_));
 sky130_fd_sc_hd__o31a_1 _12323_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A3(_05375_),
    .B1(_05163_),
    .X(_05393_));
 sky130_fd_sc_hd__xnor2_1 _12324_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__nor2_1 _12325_ (.A(_05392_),
    .B(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__and2_1 _12326_ (.A(_05392_),
    .B(_05394_),
    .X(_05396_));
 sky130_fd_sc_hd__or2_1 _12327_ (.A(_05395_),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__o21a_1 _12328_ (.A1(_05383_),
    .A2(_05385_),
    .B1(_05382_),
    .X(_05398_));
 sky130_fd_sc_hd__a21oi_1 _12329_ (.A1(_05379_),
    .A2(_05398_),
    .B1(_05387_),
    .Y(_05399_));
 sky130_fd_sc_hd__xnor2_1 _12330_ (.A(_05397_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__mux2_1 _12331_ (.A0(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_05400_),
    .S(_01249_),
    .X(_05401_));
 sky130_fd_sc_hd__and2_1 _12332_ (.A(_05290_),
    .B(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _12333_ (.A(_05402_),
    .X(_00694_));
 sky130_fd_sc_hd__inv_2 _12334_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .Y(_05403_));
 sky130_fd_sc_hd__or4_1 _12335_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .C(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .D(_05375_),
    .X(_05404_));
 sky130_fd_sc_hd__nand2_1 _12336_ (.A(_05164_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__xor2_1 _12337_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__nor2_1 _12338_ (.A(_05403_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__and2_1 _12339_ (.A(_05403_),
    .B(_05406_),
    .X(_05408_));
 sky130_fd_sc_hd__or2_1 _12340_ (.A(_05407_),
    .B(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__inv_2 _12341_ (.A(_05397_),
    .Y(_05410_));
 sky130_fd_sc_hd__a21oi_1 _12342_ (.A1(_05410_),
    .A2(_05399_),
    .B1(_05395_),
    .Y(_05411_));
 sky130_fd_sc_hd__xnor2_1 _12343_ (.A(_05409_),
    .B(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _12344_ (.A(_05142_),
    .B(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__o211a_1 _12345_ (.A1(_05140_),
    .A2(net327),
    .B1(_05141_),
    .C1(_05413_),
    .X(_00695_));
 sky130_fd_sc_hd__or2_1 _12346_ (.A(_05387_),
    .B(_05398_),
    .X(_05414_));
 sky130_fd_sc_hd__nor2_1 _12347_ (.A(_05395_),
    .B(_05407_),
    .Y(_05415_));
 sky130_fd_sc_hd__o32a_1 _12348_ (.A1(_05397_),
    .A2(_05414_),
    .A3(_05409_),
    .B1(_05415_),
    .B2(_05408_),
    .X(_05416_));
 sky130_fd_sc_hd__and2_1 _12349_ (.A(_05378_),
    .B(_05388_),
    .X(_05417_));
 sky130_fd_sc_hd__nor2_1 _12350_ (.A(_05407_),
    .B(_05408_),
    .Y(_05418_));
 sky130_fd_sc_hd__o2111ai_1 _12351_ (.A1(_05366_),
    .A2(_05370_),
    .B1(_05410_),
    .C1(_05417_),
    .D1(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__nor2_1 _12352_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05404_),
    .Y(_05420_));
 sky130_fd_sc_hd__nor2_1 _12353_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__mux2_1 _12354_ (.A0(_05421_),
    .A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .S(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_4 _12355_ (.A(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__a21o_1 _12356_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A2(_05420_),
    .B1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__xnor2_1 _12357_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__a21oi_1 _12358_ (.A1(_05416_),
    .A2(_05419_),
    .B1(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__and3_1 _12359_ (.A(_05425_),
    .B(_05416_),
    .C(_05419_),
    .X(_05427_));
 sky130_fd_sc_hd__nor2_1 _12360_ (.A(_05426_),
    .B(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__or2_1 _12361_ (.A(_05139_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(_05429_));
 sky130_fd_sc_hd__o211a_1 _12362_ (.A1(_05234_),
    .A2(_05428_),
    .B1(_05429_),
    .C1(_05343_),
    .X(_00696_));
 sky130_fd_sc_hd__buf_2 _12363_ (.A(_05423_),
    .X(_05430_));
 sky130_fd_sc_hd__and2_1 _12364_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__or2_1 _12365_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_05430_),
    .X(_05432_));
 sky130_fd_sc_hd__or2b_1 _12366_ (.A(_05431_),
    .B_N(_05432_),
    .X(_05433_));
 sky130_fd_sc_hd__a21o_1 _12367_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_05424_),
    .B1(_05426_),
    .X(_05434_));
 sky130_fd_sc_hd__xnor2_1 _12368_ (.A(_05433_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__or2_1 _12369_ (.A(_05139_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_05436_));
 sky130_fd_sc_hd__o211a_1 _12370_ (.A1(_05234_),
    .A2(_05435_),
    .B1(_05436_),
    .C1(_05343_),
    .X(_00697_));
 sky130_fd_sc_hd__or2_1 _12371_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_05430_),
    .X(_05437_));
 sky130_fd_sc_hd__nand2_1 _12372_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_05430_),
    .Y(_05438_));
 sky130_fd_sc_hd__and2_1 _12373_ (.A(_05437_),
    .B(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__o21a_1 _12374_ (.A1(_05431_),
    .A2(_05434_),
    .B1(_05432_),
    .X(_05440_));
 sky130_fd_sc_hd__nand2_1 _12375_ (.A(_05439_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__o21a_1 _12376_ (.A1(_05439_),
    .A2(_05440_),
    .B1(_01249_),
    .X(_05442_));
 sky130_fd_sc_hd__a22o_1 _12377_ (.A1(_05222_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_05441_),
    .B2(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__and2_1 _12378_ (.A(_05290_),
    .B(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_05444_),
    .X(_00698_));
 sky130_fd_sc_hd__xor2_1 _12380_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_05430_),
    .X(_05445_));
 sky130_fd_sc_hd__a21oi_1 _12381_ (.A1(_05438_),
    .A2(_05441_),
    .B1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__a31o_1 _12382_ (.A1(_05438_),
    .A2(_05441_),
    .A3(_05445_),
    .B1(_05222_),
    .X(_05447_));
 sky130_fd_sc_hd__o221a_1 _12383_ (.A1(_05142_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_05446_),
    .B2(_05447_),
    .C1(_05391_),
    .X(_00699_));
 sky130_fd_sc_hd__o31a_1 _12384_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_05423_),
    .X(_05448_));
 sky130_fd_sc_hd__a31o_1 _12385_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_05423_),
    .X(_05449_));
 sky130_fd_sc_hd__o21a_1 _12386_ (.A1(_05434_),
    .A2(_05448_),
    .B1(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__nor2_1 _12387_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05423_),
    .Y(_05451_));
 sky130_fd_sc_hd__and2_1 _12388_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05423_),
    .X(_05452_));
 sky130_fd_sc_hd__nor2_1 _12389_ (.A(_05451_),
    .B(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__xor2_1 _12390_ (.A(_05450_),
    .B(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__or2_1 _12391_ (.A(_05139_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_05455_));
 sky130_fd_sc_hd__o211a_1 _12392_ (.A1(_05234_),
    .A2(_05454_),
    .B1(_05455_),
    .C1(_05343_),
    .X(_00700_));
 sky130_fd_sc_hd__xor2_1 _12393_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_05423_),
    .X(_05456_));
 sky130_fd_sc_hd__a21oi_1 _12394_ (.A1(_05450_),
    .A2(_05453_),
    .B1(_05452_),
    .Y(_05457_));
 sky130_fd_sc_hd__nor2_1 _12395_ (.A(_05456_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__a21o_1 _12396_ (.A1(_05456_),
    .A2(_05457_),
    .B1(_05129_),
    .X(_05459_));
 sky130_fd_sc_hd__o221a_1 _12397_ (.A1(_05142_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_05458_),
    .B2(_05459_),
    .C1(_05391_),
    .X(_00701_));
 sky130_fd_sc_hd__o21a_1 _12398_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(net653),
    .B1(_05430_),
    .X(_05460_));
 sky130_fd_sc_hd__o2111a_1 _12399_ (.A1(_05434_),
    .A2(_05448_),
    .B1(_05453_),
    .C1(_05456_),
    .D1(_05449_),
    .X(_05461_));
 sky130_fd_sc_hd__or2_1 _12400_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05423_),
    .X(_05462_));
 sky130_fd_sc_hd__nand2_1 _12401_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05423_),
    .Y(_05463_));
 sky130_fd_sc_hd__and2_1 _12402_ (.A(_05462_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__o21ai_2 _12403_ (.A1(_05460_),
    .A2(_05461_),
    .B1(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__o31a_1 _12404_ (.A1(_05464_),
    .A2(_05460_),
    .A3(_05461_),
    .B1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05466_));
 sky130_fd_sc_hd__a22o_1 _12405_ (.A1(_05222_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_05465_),
    .B2(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__and2_1 _12406_ (.A(_05290_),
    .B(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__clkbuf_1 _12407_ (.A(_05468_),
    .X(_00702_));
 sky130_fd_sc_hd__xor2_1 _12408_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_05423_),
    .X(_05469_));
 sky130_fd_sc_hd__a21oi_1 _12409_ (.A1(_05463_),
    .A2(_05465_),
    .B1(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__a31o_1 _12410_ (.A1(_05463_),
    .A2(_05465_),
    .A3(_05469_),
    .B1(_05222_),
    .X(_05471_));
 sky130_fd_sc_hd__o221a_1 _12411_ (.A1(_05142_),
    .A2(net565),
    .B1(_05470_),
    .B2(_05471_),
    .C1(_05391_),
    .X(_00703_));
 sky130_fd_sc_hd__or2_1 _12412_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05430_),
    .X(_05472_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05430_),
    .Y(_05473_));
 sky130_fd_sc_hd__and2_1 _12414_ (.A(_05472_),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__o41a_1 _12415_ (.A1(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A3(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A4(net653),
    .B1(_05430_),
    .X(_05475_));
 sky130_fd_sc_hd__a31o_1 _12416_ (.A1(_05464_),
    .A2(_05461_),
    .A3(_05469_),
    .B1(_05475_),
    .X(_05476_));
 sky130_fd_sc_hd__nand2_1 _12417_ (.A(_05474_),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__o21a_1 _12418_ (.A1(_05474_),
    .A2(_05476_),
    .B1(_01249_),
    .X(_05478_));
 sky130_fd_sc_hd__a22o_1 _12419_ (.A1(_05222_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B1(_05477_),
    .B2(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__and2_1 _12420_ (.A(_05290_),
    .B(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__clkbuf_1 _12421_ (.A(_05480_),
    .X(_00704_));
 sky130_fd_sc_hd__xnor2_1 _12422_ (.A(_05275_),
    .B(_05430_),
    .Y(_05481_));
 sky130_fd_sc_hd__a21oi_1 _12423_ (.A1(_05473_),
    .A2(_05477_),
    .B1(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__a31o_1 _12424_ (.A1(_05473_),
    .A2(_05477_),
    .A3(_05481_),
    .B1(_05222_),
    .X(_05483_));
 sky130_fd_sc_hd__o221a_1 _12425_ (.A1(net536),
    .A2(_05140_),
    .B1(_05482_),
    .B2(_05483_),
    .C1(_05391_),
    .X(_00705_));
 sky130_fd_sc_hd__and2_1 _12426_ (.A(_01529_),
    .B(_02310_),
    .X(_05484_));
 sky130_fd_sc_hd__clkbuf_1 _12427_ (.A(_05484_),
    .X(_00706_));
 sky130_fd_sc_hd__inv_2 _12428_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_05485_));
 sky130_fd_sc_hd__clkbuf_4 _12429_ (.A(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__clkbuf_4 _12430_ (.A(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__clkbuf_4 _12431_ (.A(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__clkbuf_4 _12432_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05489_));
 sky130_fd_sc_hd__clkbuf_4 _12433_ (.A(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__or2_1 _12434_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__o211a_1 _12435_ (.A1(_05488_),
    .A2(net237),
    .B1(_05141_),
    .C1(_05491_),
    .X(_00707_));
 sky130_fd_sc_hd__clkbuf_4 _12436_ (.A(_05489_),
    .X(_05492_));
 sky130_fd_sc_hd__or2_1 _12437_ (.A(net207),
    .B(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__o211a_1 _12438_ (.A1(_05488_),
    .A2(net244),
    .B1(_05141_),
    .C1(_05493_),
    .X(_00708_));
 sky130_fd_sc_hd__or2_1 _12439_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B(_05492_),
    .X(_05494_));
 sky130_fd_sc_hd__o211a_1 _12440_ (.A1(_05488_),
    .A2(net149),
    .B1(_05141_),
    .C1(_05494_),
    .X(_00709_));
 sky130_fd_sc_hd__clkbuf_4 _12441_ (.A(_03619_),
    .X(_05495_));
 sky130_fd_sc_hd__or2_1 _12442_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(_05492_),
    .X(_05496_));
 sky130_fd_sc_hd__o211a_1 _12443_ (.A1(_05488_),
    .A2(net153),
    .B1(_05495_),
    .C1(_05496_),
    .X(_00710_));
 sky130_fd_sc_hd__or2_1 _12444_ (.A(net176),
    .B(_05492_),
    .X(_05497_));
 sky130_fd_sc_hd__o211a_1 _12445_ (.A1(_05488_),
    .A2(net269),
    .B1(_05495_),
    .C1(_05497_),
    .X(_00711_));
 sky130_fd_sc_hd__or2_1 _12446_ (.A(_05490_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(_05498_));
 sky130_fd_sc_hd__o211a_1 _12447_ (.A1(_05488_),
    .A2(net169),
    .B1(_05495_),
    .C1(_05498_),
    .X(_00712_));
 sky130_fd_sc_hd__clkbuf_2 _12448_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05499_));
 sky130_fd_sc_hd__clkbuf_4 _12449_ (.A(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_4 _12450_ (.A(_05489_),
    .X(_05501_));
 sky130_fd_sc_hd__nand2_1 _12451_ (.A(_05501_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .Y(_05502_));
 sky130_fd_sc_hd__o211a_1 _12452_ (.A1(_05500_),
    .A2(net350),
    .B1(_05495_),
    .C1(_05502_),
    .X(_00713_));
 sky130_fd_sc_hd__nand2_1 _12453_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .Y(_05503_));
 sky130_fd_sc_hd__or2_1 _12454_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(_05504_));
 sky130_fd_sc_hd__a21oi_1 _12455_ (.A1(_05503_),
    .A2(_05504_),
    .B1(_05203_),
    .Y(_05505_));
 sky130_fd_sc_hd__a31o_1 _12456_ (.A1(_05203_),
    .A2(_05503_),
    .A3(_05504_),
    .B1(_05487_),
    .X(_05506_));
 sky130_fd_sc_hd__o221a_1 _12457_ (.A1(_05500_),
    .A2(net552),
    .B1(_05505_),
    .B2(_05506_),
    .C1(_05391_),
    .X(_00714_));
 sky130_fd_sc_hd__and3_1 _12458_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .C(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(_05507_));
 sky130_fd_sc_hd__a21oi_1 _12459_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .Y(_05508_));
 sky130_fd_sc_hd__or2_1 _12460_ (.A(_05507_),
    .B(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__nor2_1 _12461_ (.A(_05505_),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__a21o_1 _12462_ (.A1(_05505_),
    .A2(_05509_),
    .B1(_05487_),
    .X(_05511_));
 sky130_fd_sc_hd__o221a_1 _12463_ (.A1(_05500_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B1(_05510_),
    .B2(_05511_),
    .C1(_05391_),
    .X(_00715_));
 sky130_fd_sc_hd__nand2_1 _12464_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05507_),
    .Y(_05512_));
 sky130_fd_sc_hd__o31a_1 _12465_ (.A1(_05203_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A3(_05504_),
    .B1(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__and2_1 _12466_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__o21ai_1 _12467_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(_05513_),
    .B1(_05501_),
    .Y(_05515_));
 sky130_fd_sc_hd__o221a_1 _12468_ (.A1(_05500_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B1(_05514_),
    .B2(_05515_),
    .C1(_05391_),
    .X(_00716_));
 sky130_fd_sc_hd__or3_1 _12469_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .C(_05504_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_1 _12470_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_05507_),
    .Y(_05517_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(_05516_),
    .A1(_05517_),
    .S(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05518_));
 sky130_fd_sc_hd__and2_1 _12472_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__o21ai_1 _12473_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_05518_),
    .B1(_05490_),
    .Y(_05520_));
 sky130_fd_sc_hd__o221a_1 _12474_ (.A1(_05500_),
    .A2(net519),
    .B1(_05519_),
    .B2(_05520_),
    .C1(_05391_),
    .X(_00717_));
 sky130_fd_sc_hd__clkbuf_4 _12475_ (.A(_05489_),
    .X(_05521_));
 sky130_fd_sc_hd__or3_1 _12476_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(_05516_),
    .X(_05522_));
 sky130_fd_sc_hd__o21ai_1 _12477_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_05516_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_05523_));
 sky130_fd_sc_hd__a21oi_1 _12478_ (.A1(_05522_),
    .A2(_05523_),
    .B1(_05203_),
    .Y(_05524_));
 sky130_fd_sc_hd__inv_2 _12479_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_05525_));
 sky130_fd_sc_hd__clkbuf_4 _12480_ (.A(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__a31oi_1 _12481_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A3(_05507_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_05527_));
 sky130_fd_sc_hd__and4_1 _12482_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .D(_05507_),
    .X(_05528_));
 sky130_fd_sc_hd__o31ai_1 _12483_ (.A1(_05526_),
    .A2(_05527_),
    .A3(_05528_),
    .B1(_05490_),
    .Y(_05529_));
 sky130_fd_sc_hd__o221a_1 _12484_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B1(_05524_),
    .B2(_05529_),
    .C1(_05391_),
    .X(_00718_));
 sky130_fd_sc_hd__inv_2 _12485_ (.A(_05522_),
    .Y(_05530_));
 sky130_fd_sc_hd__mux2_1 _12486_ (.A0(_05530_),
    .A1(_05528_),
    .S(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05531_));
 sky130_fd_sc_hd__xnor2_1 _12487_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(_05501_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__o211a_1 _12489_ (.A1(_05500_),
    .A2(net584),
    .B1(_05495_),
    .C1(_05533_),
    .X(_00719_));
 sky130_fd_sc_hd__nand2_1 _12490_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_05528_),
    .Y(_05534_));
 sky130_fd_sc_hd__or2_1 _12491_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_05522_),
    .X(_05535_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(_05534_),
    .A1(_05535_),
    .S(_05526_),
    .X(_05536_));
 sky130_fd_sc_hd__o21ai_1 _12493_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_05536_),
    .B1(_05489_),
    .Y(_05537_));
 sky130_fd_sc_hd__a21o_1 _12494_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_05536_),
    .B1(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__o211a_1 _12495_ (.A1(_05500_),
    .A2(net602),
    .B1(_05495_),
    .C1(_05538_),
    .X(_00720_));
 sky130_fd_sc_hd__and3_1 _12496_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_05528_),
    .X(_05539_));
 sky130_fd_sc_hd__nand2_1 _12497_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__o31a_1 _12498_ (.A1(_05203_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(_05535_),
    .B1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__and2_1 _12499_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__o21ai_1 _12500_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_05541_),
    .B1(_05490_),
    .Y(_05543_));
 sky130_fd_sc_hd__clkbuf_4 _12501_ (.A(_04538_),
    .X(_05544_));
 sky130_fd_sc_hd__o221a_1 _12502_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_05542_),
    .B2(_05543_),
    .C1(_05544_),
    .X(_00721_));
 sky130_fd_sc_hd__nand3_1 _12503_ (.A(_05203_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C(_05539_),
    .Y(_05545_));
 sky130_fd_sc_hd__o41a_1 _12504_ (.A1(_05203_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A3(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A4(_05535_),
    .B1(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__nor2_1 _12505_ (.A(net529),
    .B(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__a21o_1 _12506_ (.A1(net615),
    .A2(_05546_),
    .B1(_05487_),
    .X(_05548_));
 sky130_fd_sc_hd__o221a_1 _12507_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_05547_),
    .B2(_05548_),
    .C1(_05544_),
    .X(_00722_));
 sky130_fd_sc_hd__or4_1 _12508_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .D(_05535_),
    .X(_05549_));
 sky130_fd_sc_hd__and3_1 _12509_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .C(_05539_),
    .X(_05550_));
 sky130_fd_sc_hd__nand2_1 _12510_ (.A(_05203_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__o21a_1 _12511_ (.A1(_05203_),
    .A2(_05549_),
    .B1(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__and2_1 _12512_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__o21ai_1 _12513_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_05552_),
    .B1(_05490_),
    .Y(_05554_));
 sky130_fd_sc_hd__o221a_1 _12514_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_05553_),
    .B2(_05554_),
    .C1(_05544_),
    .X(_00723_));
 sky130_fd_sc_hd__nand2_1 _12515_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_05550_),
    .Y(_05555_));
 sky130_fd_sc_hd__or2_1 _12516_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_05549_),
    .X(_05556_));
 sky130_fd_sc_hd__mux2_1 _12517_ (.A0(_05555_),
    .A1(_05556_),
    .S(_05526_),
    .X(_05557_));
 sky130_fd_sc_hd__nor2_1 _12518_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__a21o_1 _12519_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05557_),
    .B1(_05487_),
    .X(_05559_));
 sky130_fd_sc_hd__o221a_1 _12520_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_05558_),
    .B2(_05559_),
    .C1(_05544_),
    .X(_00724_));
 sky130_fd_sc_hd__o21a_1 _12521_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05556_),
    .B1(_05526_),
    .X(_05560_));
 sky130_fd_sc_hd__a31o_1 _12522_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_05550_),
    .B1(_05526_),
    .X(_05561_));
 sky130_fd_sc_hd__or2b_1 _12523_ (.A(_05560_),
    .B_N(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__xnor2_1 _12524_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__or2_1 _12525_ (.A(_05492_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_05564_));
 sky130_fd_sc_hd__o211a_1 _12526_ (.A1(_05488_),
    .A2(_05563_),
    .B1(_05564_),
    .C1(_05343_),
    .X(_00725_));
 sky130_fd_sc_hd__a21oi_1 _12527_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_05561_),
    .B1(_05560_),
    .Y(_05565_));
 sky130_fd_sc_hd__clkbuf_4 _12528_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05566_));
 sky130_fd_sc_hd__buf_2 _12529_ (.A(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__or2_1 _12530_ (.A(_05492_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__o211a_1 _12531_ (.A1(_05488_),
    .A2(_05565_),
    .B1(_05568_),
    .C1(_05343_),
    .X(_00726_));
 sky130_fd_sc_hd__inv_2 _12532_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .Y(_05569_));
 sky130_fd_sc_hd__nor2_1 _12533_ (.A(_05569_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_05570_));
 sky130_fd_sc_hd__a21o_1 _12534_ (.A1(_05569_),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_05487_),
    .X(_05571_));
 sky130_fd_sc_hd__o221a_1 _12535_ (.A1(_05521_),
    .A2(net471),
    .B1(_05570_),
    .B2(_05571_),
    .C1(_05544_),
    .X(_00727_));
 sky130_fd_sc_hd__and2b_1 _12536_ (.A_N(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .X(_05572_));
 sky130_fd_sc_hd__xnor2_1 _12537_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__xnor2_1 _12538_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__xor2_1 _12539_ (.A(_05570_),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__or2_1 _12540_ (.A(_05492_),
    .B(net607),
    .X(_05576_));
 sky130_fd_sc_hd__o211a_1 _12541_ (.A1(_05488_),
    .A2(_05575_),
    .B1(_05576_),
    .C1(_05343_),
    .X(_00728_));
 sky130_fd_sc_hd__o21a_1 _12542_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_05525_),
    .X(_05577_));
 sky130_fd_sc_hd__xnor2_1 _12543_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__nor2_1 _12544_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand2_1 _12545_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_05578_),
    .Y(_05580_));
 sky130_fd_sc_hd__or2b_1 _12546_ (.A(_05579_),
    .B_N(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__nand2_1 _12547_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_05573_),
    .Y(_05582_));
 sky130_fd_sc_hd__o21a_1 _12548_ (.A1(_05570_),
    .A2(_05574_),
    .B1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__a21o_1 _12549_ (.A1(_05581_),
    .A2(_05583_),
    .B1(_05485_),
    .X(_05584_));
 sky130_fd_sc_hd__nor2_1 _12550_ (.A(_05581_),
    .B(_05583_),
    .Y(_05585_));
 sky130_fd_sc_hd__a2bb2o_1 _12551_ (.A1_N(_05584_),
    .A2_N(_05585_),
    .B1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B2(_05486_),
    .X(_05586_));
 sky130_fd_sc_hd__and2_1 _12552_ (.A(_05290_),
    .B(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__clkbuf_1 _12553_ (.A(_05587_),
    .X(_00729_));
 sky130_fd_sc_hd__o31a_1 _12554_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A3(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_05526_),
    .X(_05588_));
 sky130_fd_sc_hd__xnor2_1 _12555_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__and2_1 _12556_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__or2_1 _12557_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_05589_),
    .X(_05591_));
 sky130_fd_sc_hd__and2b_1 _12558_ (.A_N(_05590_),
    .B(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__o21ai_1 _12559_ (.A1(_05579_),
    .A2(_05583_),
    .B1(_05580_),
    .Y(_05593_));
 sky130_fd_sc_hd__xor2_1 _12560_ (.A(_05592_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_05594_),
    .S(_05489_),
    .X(_05595_));
 sky130_fd_sc_hd__and2_1 _12562_ (.A(_05290_),
    .B(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_1 _12563_ (.A(_05596_),
    .X(_00730_));
 sky130_fd_sc_hd__a21o_1 _12564_ (.A1(_05591_),
    .A2(_05593_),
    .B1(_05590_),
    .X(_05597_));
 sky130_fd_sc_hd__or4_2 _12565_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .C(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .D(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .X(_05598_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(_05526_),
    .B(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__xor2_1 _12567_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__and2_1 _12568_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__nor2_1 _12569_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_05600_),
    .Y(_05602_));
 sky130_fd_sc_hd__nor2_1 _12570_ (.A(_05601_),
    .B(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__xor2_1 _12571_ (.A(_05597_),
    .B(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__or2_1 _12572_ (.A(_05492_),
    .B(net498),
    .X(_05605_));
 sky130_fd_sc_hd__o211a_1 _12573_ (.A1(_05488_),
    .A2(_05604_),
    .B1(_05605_),
    .C1(_05343_),
    .X(_00731_));
 sky130_fd_sc_hd__o21a_1 _12574_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(_05598_),
    .B1(_05526_),
    .X(_05606_));
 sky130_fd_sc_hd__xnor2_1 _12575_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__nand2_2 _12576_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__or2_1 _12577_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_05607_),
    .X(_05609_));
 sky130_fd_sc_hd__nand2_1 _12578_ (.A(_05608_),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__a21o_1 _12579_ (.A1(_05597_),
    .A2(_05603_),
    .B1(_05601_),
    .X(_05611_));
 sky130_fd_sc_hd__and2_1 _12580_ (.A(_05610_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__o21ai_1 _12581_ (.A1(_05610_),
    .A2(_05611_),
    .B1(_05490_),
    .Y(_05613_));
 sky130_fd_sc_hd__o221a_1 _12582_ (.A1(_05521_),
    .A2(net352),
    .B1(_05612_),
    .B2(_05613_),
    .C1(_05544_),
    .X(_00732_));
 sky130_fd_sc_hd__inv_2 _12583_ (.A(net586),
    .Y(_05614_));
 sky130_fd_sc_hd__nor2_1 _12584_ (.A(_05501_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_1 _12585_ (.A(_05609_),
    .B(_05611_),
    .Y(_05616_));
 sky130_fd_sc_hd__o31a_1 _12586_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A3(_05598_),
    .B1(_05526_),
    .X(_05617_));
 sky130_fd_sc_hd__xnor2_1 _12587_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _12588_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _12589_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_1 _12590_ (.A(_05619_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__a31o_1 _12591_ (.A1(_05608_),
    .A2(_05616_),
    .A3(_05621_),
    .B1(_05486_),
    .X(_05622_));
 sky130_fd_sc_hd__a21o_1 _12592_ (.A1(_05608_),
    .A2(_05616_),
    .B1(_05621_),
    .X(_05623_));
 sky130_fd_sc_hd__and2b_1 _12593_ (.A_N(_05622_),
    .B(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__o21a_1 _12594_ (.A1(_05615_),
    .A2(_05624_),
    .B1(_04961_),
    .X(_00733_));
 sky130_fd_sc_hd__o41a_1 _12595_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A3(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A4(_05598_),
    .B1(_05525_),
    .X(_05625_));
 sky130_fd_sc_hd__xnor2_1 _12596_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__and2_1 _12597_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__nor2_1 _12598_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_05626_),
    .Y(_05628_));
 sky130_fd_sc_hd__nor2_1 _12599_ (.A(_05627_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__a21oi_1 _12600_ (.A1(_05619_),
    .A2(_05623_),
    .B1(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__a31o_1 _12601_ (.A1(_05619_),
    .A2(_05623_),
    .A3(_05629_),
    .B1(_05487_),
    .X(_05631_));
 sky130_fd_sc_hd__o221a_1 _12602_ (.A1(_05521_),
    .A2(net399),
    .B1(_05630_),
    .B2(_05631_),
    .C1(_05544_),
    .X(_00734_));
 sky130_fd_sc_hd__buf_2 _12603_ (.A(_05487_),
    .X(_05632_));
 sky130_fd_sc_hd__inv_2 _12604_ (.A(_05608_),
    .Y(_05633_));
 sky130_fd_sc_hd__o211ai_1 _12605_ (.A1(_05601_),
    .A2(_05633_),
    .B1(_05609_),
    .C1(_05629_),
    .Y(_05634_));
 sky130_fd_sc_hd__inv_2 _12606_ (.A(_05627_),
    .Y(_05635_));
 sky130_fd_sc_hd__o221a_1 _12607_ (.A1(_05619_),
    .A2(_05628_),
    .B1(_05634_),
    .B2(_05621_),
    .C1(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__nand3_1 _12608_ (.A(_05603_),
    .B(_05608_),
    .C(_05609_),
    .Y(_05637_));
 sky130_fd_sc_hd__or4bb_1 _12609_ (.A(_05621_),
    .B(_05637_),
    .C_N(_05629_),
    .D_N(_05597_),
    .X(_05638_));
 sky130_fd_sc_hd__nor2_1 _12610_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05625_),
    .Y(_05639_));
 sky130_fd_sc_hd__a21o_1 _12611_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_05526_),
    .B1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__clkbuf_4 _12612_ (.A(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__xnor2_1 _12613_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__a21oi_1 _12614_ (.A1(_05636_),
    .A2(_05638_),
    .B1(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__and3_1 _12615_ (.A(_05642_),
    .B(_05636_),
    .C(_05638_),
    .X(_05644_));
 sky130_fd_sc_hd__nor2_1 _12616_ (.A(_05643_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__or2_1 _12617_ (.A(_05492_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_05646_));
 sky130_fd_sc_hd__o211a_1 _12618_ (.A1(_05632_),
    .A2(_05645_),
    .B1(_05646_),
    .C1(_05343_),
    .X(_00735_));
 sky130_fd_sc_hd__xor2_1 _12619_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_05641_),
    .X(_05647_));
 sky130_fd_sc_hd__buf_2 _12620_ (.A(_05641_),
    .X(_05648_));
 sky130_fd_sc_hd__a21o_1 _12621_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_05648_),
    .B1(_05643_),
    .X(_05649_));
 sky130_fd_sc_hd__xor2_1 _12622_ (.A(_05647_),
    .B(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__or2_1 _12623_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_05651_));
 sky130_fd_sc_hd__o211a_1 _12624_ (.A1(_05632_),
    .A2(_05650_),
    .B1(_05651_),
    .C1(_05343_),
    .X(_00736_));
 sky130_fd_sc_hd__buf_2 _12625_ (.A(_01252_),
    .X(_05652_));
 sky130_fd_sc_hd__o21a_1 _12626_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_05648_),
    .X(_05653_));
 sky130_fd_sc_hd__o21a_1 _12627_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_05648_),
    .B1(_05643_),
    .X(_05654_));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_05641_),
    .Y(_05655_));
 sky130_fd_sc_hd__or2_1 _12629_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_05640_),
    .X(_05656_));
 sky130_fd_sc_hd__and2_1 _12630_ (.A(_05655_),
    .B(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__o21ai_2 _12631_ (.A1(_05653_),
    .A2(_05654_),
    .B1(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__or3_1 _12632_ (.A(_05657_),
    .B(_05653_),
    .C(_05654_),
    .X(_05659_));
 sky130_fd_sc_hd__and2_1 _12633_ (.A(_05485_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_05660_));
 sky130_fd_sc_hd__a31o_1 _12634_ (.A1(_05489_),
    .A2(_05658_),
    .A3(_05659_),
    .B1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__and2_1 _12635_ (.A(_05652_),
    .B(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _12636_ (.A(_05662_),
    .X(_00737_));
 sky130_fd_sc_hd__xor2_2 _12637_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_05641_),
    .X(_05663_));
 sky130_fd_sc_hd__a21oi_1 _12638_ (.A1(_05655_),
    .A2(_05658_),
    .B1(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__a31o_1 _12639_ (.A1(_05655_),
    .A2(_05658_),
    .A3(_05663_),
    .B1(_05487_),
    .X(_05665_));
 sky130_fd_sc_hd__o221a_1 _12640_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_05664_),
    .B2(_05665_),
    .C1(_05544_),
    .X(_00738_));
 sky130_fd_sc_hd__nand2_1 _12641_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05641_),
    .Y(_05666_));
 sky130_fd_sc_hd__or2_1 _12642_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05641_),
    .X(_05667_));
 sky130_fd_sc_hd__and2_1 _12643_ (.A(_05666_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__and4_1 _12644_ (.A(_05643_),
    .B(_05647_),
    .C(_05657_),
    .D(_05663_),
    .X(_05669_));
 sky130_fd_sc_hd__o41a_2 _12645_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A3(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A4(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_05648_),
    .X(_05670_));
 sky130_fd_sc_hd__or3_1 _12646_ (.A(_05668_),
    .B(_05669_),
    .C(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__o21ai_1 _12647_ (.A1(_05669_),
    .A2(_05670_),
    .B1(_05668_),
    .Y(_05672_));
 sky130_fd_sc_hd__and2_1 _12648_ (.A(_05671_),
    .B(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__or2_1 _12649_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_05674_));
 sky130_fd_sc_hd__buf_4 _12650_ (.A(_04455_),
    .X(_05675_));
 sky130_fd_sc_hd__o211a_1 _12651_ (.A1(_05632_),
    .A2(_05673_),
    .B1(_05674_),
    .C1(_05675_),
    .X(_00739_));
 sky130_fd_sc_hd__xor2_1 _12652_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_05641_),
    .X(_05676_));
 sky130_fd_sc_hd__a21oi_1 _12653_ (.A1(_05666_),
    .A2(_05672_),
    .B1(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__a31o_1 _12654_ (.A1(_05666_),
    .A2(_05672_),
    .A3(_05676_),
    .B1(_05486_),
    .X(_05678_));
 sky130_fd_sc_hd__o221a_1 _12655_ (.A1(_05521_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_05677_),
    .B2(_05678_),
    .C1(_05544_),
    .X(_00740_));
 sky130_fd_sc_hd__and2_1 _12656_ (.A(_05487_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .X(_05679_));
 sky130_fd_sc_hd__o21a_1 _12657_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_05648_),
    .X(_05680_));
 sky130_fd_sc_hd__and2_1 _12658_ (.A(_05668_),
    .B(_05676_),
    .X(_05681_));
 sky130_fd_sc_hd__o21a_1 _12659_ (.A1(_05669_),
    .A2(_05670_),
    .B1(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__xor2_1 _12660_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_05641_),
    .X(_05683_));
 sky130_fd_sc_hd__o21a_1 _12661_ (.A1(_05680_),
    .A2(_05682_),
    .B1(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__or3_1 _12662_ (.A(_05683_),
    .B(_05680_),
    .C(_05682_),
    .X(_05685_));
 sky130_fd_sc_hd__and3b_1 _12663_ (.A_N(_05684_),
    .B(_05685_),
    .C(_05492_),
    .X(_05686_));
 sky130_fd_sc_hd__o21a_1 _12664_ (.A1(_05679_),
    .A2(_05686_),
    .B1(_04961_),
    .X(_00741_));
 sky130_fd_sc_hd__a21o_1 _12665_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_05648_),
    .B1(_05684_),
    .X(_05687_));
 sky130_fd_sc_hd__xor2_1 _12666_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_05641_),
    .X(_05688_));
 sky130_fd_sc_hd__xor2_1 _12667_ (.A(_05687_),
    .B(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__or2_1 _12668_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(_05690_));
 sky130_fd_sc_hd__o211a_1 _12669_ (.A1(_05632_),
    .A2(_05689_),
    .B1(_05690_),
    .C1(_05675_),
    .X(_00742_));
 sky130_fd_sc_hd__and4_1 _12670_ (.A(_05669_),
    .B(_05683_),
    .C(_05681_),
    .D(_05688_),
    .X(_05691_));
 sky130_fd_sc_hd__o41a_1 _12671_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A3(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A4(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_05648_),
    .X(_05692_));
 sky130_fd_sc_hd__or2_1 _12672_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05648_),
    .X(_05693_));
 sky130_fd_sc_hd__nand2_1 _12673_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05648_),
    .Y(_05694_));
 sky130_fd_sc_hd__and2_1 _12674_ (.A(_05693_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__o31ai_2 _12675_ (.A1(_05670_),
    .A2(_05691_),
    .A3(_05692_),
    .B1(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__o41a_1 _12676_ (.A1(_05670_),
    .A2(_05695_),
    .A3(_05691_),
    .A4(_05692_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05697_));
 sky130_fd_sc_hd__a22o_1 _12677_ (.A1(_05486_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B1(_05696_),
    .B2(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__and2_1 _12678_ (.A(_05652_),
    .B(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_1 _12679_ (.A(_05699_),
    .X(_00743_));
 sky130_fd_sc_hd__xor2_1 _12680_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_05648_),
    .X(_05700_));
 sky130_fd_sc_hd__a21oi_1 _12681_ (.A1(_05694_),
    .A2(_05696_),
    .B1(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__a31o_1 _12682_ (.A1(_05694_),
    .A2(_05696_),
    .A3(_05700_),
    .B1(_05486_),
    .X(_05702_));
 sky130_fd_sc_hd__o221a_1 _12683_ (.A1(_05501_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B1(_05701_),
    .B2(_05702_),
    .C1(_05544_),
    .X(_00744_));
 sky130_fd_sc_hd__and2_1 _12684_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_05703_));
 sky130_fd_sc_hd__nor2_1 _12685_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ai_1 _12686_ (.A1(_05703_),
    .A2(_05704_),
    .B1(_05501_),
    .Y(_05705_));
 sky130_fd_sc_hd__o211a_1 _12687_ (.A1(_05500_),
    .A2(net315),
    .B1(_05495_),
    .C1(_05705_),
    .X(_00745_));
 sky130_fd_sc_hd__and2b_1 _12688_ (.A_N(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_05706_));
 sky130_fd_sc_hd__xnor2_1 _12689_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__xnor2_1 _12690_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__xor2_1 _12691_ (.A(_05703_),
    .B(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__or2_1 _12692_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_05710_));
 sky130_fd_sc_hd__o211a_1 _12693_ (.A1(_05632_),
    .A2(_05709_),
    .B1(_05710_),
    .C1(_05675_),
    .X(_00746_));
 sky130_fd_sc_hd__o21a_1 _12694_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_05525_),
    .X(_05711_));
 sky130_fd_sc_hd__xnor2_1 _12695_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__and2_1 _12696_ (.A(_05359_),
    .B(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__nor2_1 _12697_ (.A(_05359_),
    .B(_05712_),
    .Y(_05714_));
 sky130_fd_sc_hd__nor2_1 _12698_ (.A(_05713_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__and2b_1 _12699_ (.A_N(_05707_),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_05716_));
 sky130_fd_sc_hd__a21o_1 _12700_ (.A1(_05703_),
    .A2(_05708_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(_05715_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__o21a_1 _12702_ (.A1(_05715_),
    .A2(_05717_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05719_));
 sky130_fd_sc_hd__a22o_1 _12703_ (.A1(_05486_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_05718_),
    .B2(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__and2_1 _12704_ (.A(_05652_),
    .B(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__clkbuf_1 _12705_ (.A(_05721_),
    .X(_00747_));
 sky130_fd_sc_hd__a21o_1 _12706_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_05525_),
    .B1(_05711_),
    .X(_05722_));
 sky130_fd_sc_hd__xor2_1 _12707_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__and2_1 _12708_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__or2_1 _12709_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_05723_),
    .X(_05725_));
 sky130_fd_sc_hd__or2b_1 _12710_ (.A(_05724_),
    .B_N(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _12711_ (.A(_05359_),
    .B(_05712_),
    .Y(_05727_));
 sky130_fd_sc_hd__a21o_1 _12712_ (.A1(_05727_),
    .A2(_05717_),
    .B1(_05714_),
    .X(_05728_));
 sky130_fd_sc_hd__xnor2_1 _12713_ (.A(_05726_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A1(_05729_),
    .S(_05489_),
    .X(_05730_));
 sky130_fd_sc_hd__and2_1 _12715_ (.A(_05652_),
    .B(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_1 _12716_ (.A(_05731_),
    .X(_00748_));
 sky130_fd_sc_hd__a21oi_2 _12717_ (.A1(_05725_),
    .A2(_05728_),
    .B1(_05724_),
    .Y(_05732_));
 sky130_fd_sc_hd__inv_2 _12718_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_05733_));
 sky130_fd_sc_hd__or4_2 _12719_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .C(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .D(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_1 _12720_ (.A(_05525_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__xor2_1 _12721_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__nor2_1 _12722_ (.A(_05733_),
    .B(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__and2_1 _12723_ (.A(_05733_),
    .B(_05736_),
    .X(_05738_));
 sky130_fd_sc_hd__or2_1 _12724_ (.A(_05737_),
    .B(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__nor2_1 _12725_ (.A(_05732_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__and2_1 _12726_ (.A(_05732_),
    .B(_05739_),
    .X(_05741_));
 sky130_fd_sc_hd__nor2_1 _12727_ (.A(_05740_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__or2_1 _12728_ (.A(_05499_),
    .B(net641),
    .X(_05743_));
 sky130_fd_sc_hd__o211a_1 _12729_ (.A1(_05632_),
    .A2(_05742_),
    .B1(_05743_),
    .C1(_05675_),
    .X(_00749_));
 sky130_fd_sc_hd__o21a_1 _12730_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_05734_),
    .B1(_05525_),
    .X(_05744_));
 sky130_fd_sc_hd__xor2_1 _12731_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__and2_1 _12732_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__or2_1 _12733_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_05745_),
    .X(_05747_));
 sky130_fd_sc_hd__or2b_1 _12734_ (.A(_05746_),
    .B_N(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__o21a_1 _12735_ (.A1(_05737_),
    .A2(_05740_),
    .B1(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__o31ai_1 _12736_ (.A1(_05737_),
    .A2(_05740_),
    .A3(_05748_),
    .B1(_05490_),
    .Y(_05750_));
 sky130_fd_sc_hd__buf_4 _12737_ (.A(_04538_),
    .X(_05751_));
 sky130_fd_sc_hd__o221a_1 _12738_ (.A1(_05501_),
    .A2(net311),
    .B1(_05749_),
    .B2(_05750_),
    .C1(_05751_),
    .X(_00750_));
 sky130_fd_sc_hd__or2_1 _12739_ (.A(_05739_),
    .B(_05748_),
    .X(_05752_));
 sky130_fd_sc_hd__or2_1 _12740_ (.A(_05732_),
    .B(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__o21ai_2 _12741_ (.A1(_05737_),
    .A2(_05746_),
    .B1(_05747_),
    .Y(_05754_));
 sky130_fd_sc_hd__inv_2 _12742_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .Y(_05755_));
 sky130_fd_sc_hd__or3_1 _12743_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .C(_05734_),
    .X(_05756_));
 sky130_fd_sc_hd__and2_1 _12744_ (.A(_05525_),
    .B(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__xnor2_1 _12745_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__nor2_1 _12746_ (.A(_05755_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__and2_1 _12747_ (.A(_05755_),
    .B(_05758_),
    .X(_05760_));
 sky130_fd_sc_hd__or2_1 _12748_ (.A(_05759_),
    .B(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__a21o_1 _12749_ (.A1(_05753_),
    .A2(_05754_),
    .B1(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__o211a_1 _12750_ (.A1(_05732_),
    .A2(_05752_),
    .B1(_05754_),
    .C1(_05761_),
    .X(_05763_));
 sky130_fd_sc_hd__nor2_1 _12751_ (.A(_05485_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__a22o_1 _12752_ (.A1(_05486_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1(_05762_),
    .B2(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__and2_1 _12753_ (.A(_05652_),
    .B(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__clkbuf_1 _12754_ (.A(_05766_),
    .X(_00751_));
 sky130_fd_sc_hd__nor2_1 _12755_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_05756_),
    .Y(_05767_));
 sky130_fd_sc_hd__and2_1 _12756_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__or2_1 _12757_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05769_));
 sky130_fd_sc_hd__nand2_1 _12758_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_05770_));
 sky130_fd_sc_hd__o21ai_1 _12759_ (.A1(_05767_),
    .A2(_05769_),
    .B1(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21a_1 _12760_ (.A1(_05768_),
    .A2(_05771_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_05772_));
 sky130_fd_sc_hd__nor3_1 _12761_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_05768_),
    .C(_05771_),
    .Y(_05773_));
 sky130_fd_sc_hd__or2_1 _12762_ (.A(_05772_),
    .B(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__or2b_1 _12763_ (.A(_05759_),
    .B_N(_05762_),
    .X(_05775_));
 sky130_fd_sc_hd__o21ai_1 _12764_ (.A1(_05774_),
    .A2(_05775_),
    .B1(_05489_),
    .Y(_05776_));
 sky130_fd_sc_hd__a21o_1 _12765_ (.A1(_05774_),
    .A2(_05775_),
    .B1(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__o211a_1 _12766_ (.A1(_05500_),
    .A2(net264),
    .B1(_05495_),
    .C1(_05777_),
    .X(_00752_));
 sky130_fd_sc_hd__nor2_1 _12767_ (.A(_05759_),
    .B(_05772_),
    .Y(_05778_));
 sky130_fd_sc_hd__o32a_1 _12768_ (.A1(_05761_),
    .A2(_05754_),
    .A3(_05774_),
    .B1(_05778_),
    .B2(_05773_),
    .X(_05779_));
 sky130_fd_sc_hd__or4_1 _12769_ (.A(_05732_),
    .B(_05761_),
    .C(_05752_),
    .D(_05774_),
    .X(_05780_));
 sky130_fd_sc_hd__clkbuf_4 _12770_ (.A(_05771_),
    .X(_05781_));
 sky130_fd_sc_hd__xnor2_1 _12771_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__a21oi_1 _12772_ (.A1(_05779_),
    .A2(_05780_),
    .B1(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__and3_1 _12773_ (.A(_05782_),
    .B(_05779_),
    .C(_05780_),
    .X(_05784_));
 sky130_fd_sc_hd__o21ai_1 _12774_ (.A1(_05783_),
    .A2(_05784_),
    .B1(_05501_),
    .Y(_05785_));
 sky130_fd_sc_hd__o211a_1 _12775_ (.A1(_05500_),
    .A2(net634),
    .B1(_05495_),
    .C1(_05785_),
    .X(_00753_));
 sky130_fd_sc_hd__nor2_1 _12776_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_05781_),
    .Y(_05786_));
 sky130_fd_sc_hd__and2_1 _12777_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_05781_),
    .X(_05787_));
 sky130_fd_sc_hd__nor2_1 _12778_ (.A(_05786_),
    .B(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__clkbuf_4 _12779_ (.A(_05781_),
    .X(_05789_));
 sky130_fd_sc_hd__a21oi_1 _12780_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_05789_),
    .B1(_05783_),
    .Y(_05790_));
 sky130_fd_sc_hd__xnor2_1 _12781_ (.A(_05788_),
    .B(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__or2_1 _12782_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_05792_));
 sky130_fd_sc_hd__o211a_1 _12783_ (.A1(_05632_),
    .A2(_05791_),
    .B1(_05792_),
    .C1(_05675_),
    .X(_00754_));
 sky130_fd_sc_hd__nor2_1 _12784_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_05781_),
    .Y(_05793_));
 sky130_fd_sc_hd__and2_1 _12785_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_05781_),
    .X(_05794_));
 sky130_fd_sc_hd__nor2_1 _12786_ (.A(_05793_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__o21bai_1 _12787_ (.A1(_05786_),
    .A2(_05790_),
    .B1_N(_05787_),
    .Y(_05796_));
 sky130_fd_sc_hd__xor2_1 _12788_ (.A(_05795_),
    .B(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__mux2_1 _12789_ (.A0(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A1(_05797_),
    .S(_05489_),
    .X(_05798_));
 sky130_fd_sc_hd__and2_1 _12790_ (.A(_05652_),
    .B(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_1 _12791_ (.A(_05799_),
    .X(_00755_));
 sky130_fd_sc_hd__a21oi_1 _12792_ (.A1(_05795_),
    .A2(_05796_),
    .B1(_05794_),
    .Y(_05800_));
 sky130_fd_sc_hd__xor2_1 _12793_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_05781_),
    .X(_05801_));
 sky130_fd_sc_hd__and2_1 _12794_ (.A(_05800_),
    .B(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__o21ai_1 _12795_ (.A1(_05800_),
    .A2(_05801_),
    .B1(_05490_),
    .Y(_05803_));
 sky130_fd_sc_hd__o221a_1 _12796_ (.A1(_05501_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_05802_),
    .B2(_05803_),
    .C1(_05751_),
    .X(_00756_));
 sky130_fd_sc_hd__nor2_1 _12797_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05781_),
    .Y(_05804_));
 sky130_fd_sc_hd__and2_1 _12798_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05781_),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _12799_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__and4_1 _12800_ (.A(_05783_),
    .B(_05788_),
    .C(_05795_),
    .D(_05801_),
    .X(_05807_));
 sky130_fd_sc_hd__o41a_1 _12801_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A4(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_05789_),
    .X(_05808_));
 sky130_fd_sc_hd__or2_1 _12802_ (.A(_05807_),
    .B(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__xor2_1 _12803_ (.A(_05806_),
    .B(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__or2_1 _12804_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_05811_));
 sky130_fd_sc_hd__o211a_1 _12805_ (.A1(_05632_),
    .A2(_05810_),
    .B1(_05811_),
    .C1(_05675_),
    .X(_00757_));
 sky130_fd_sc_hd__xor2_1 _12806_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_05781_),
    .X(_05812_));
 sky130_fd_sc_hd__a21o_1 _12807_ (.A1(_05806_),
    .A2(_05809_),
    .B1(_05805_),
    .X(_05813_));
 sky130_fd_sc_hd__xor2_1 _12808_ (.A(_05812_),
    .B(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__or2_1 _12809_ (.A(_05499_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_05815_));
 sky130_fd_sc_hd__o211a_1 _12810_ (.A1(_05632_),
    .A2(_05814_),
    .B1(_05815_),
    .C1(_05675_),
    .X(_00758_));
 sky130_fd_sc_hd__o21a_1 _12811_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_05789_),
    .X(_05816_));
 sky130_fd_sc_hd__and2_1 _12812_ (.A(_05806_),
    .B(_05812_),
    .X(_05817_));
 sky130_fd_sc_hd__and2_1 _12813_ (.A(_05809_),
    .B(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__or2_1 _12814_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05789_),
    .X(_05819_));
 sky130_fd_sc_hd__nand2_1 _12815_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05789_),
    .Y(_05820_));
 sky130_fd_sc_hd__and2_1 _12816_ (.A(_05819_),
    .B(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__o21ai_1 _12817_ (.A1(_05816_),
    .A2(_05818_),
    .B1(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__o31a_1 _12818_ (.A1(_05821_),
    .A2(_05816_),
    .A3(_05818_),
    .B1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05823_));
 sky130_fd_sc_hd__a22o_1 _12819_ (.A1(_05486_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_05822_),
    .B2(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__and2_1 _12820_ (.A(_05652_),
    .B(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_1 _12821_ (.A(_05825_),
    .X(_00759_));
 sky130_fd_sc_hd__xor2_2 _12822_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_05789_),
    .X(_05826_));
 sky130_fd_sc_hd__a21oi_1 _12823_ (.A1(_05820_),
    .A2(_05822_),
    .B1(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__a31o_1 _12824_ (.A1(_05820_),
    .A2(_05822_),
    .A3(_05826_),
    .B1(_05486_),
    .X(_05828_));
 sky130_fd_sc_hd__o221a_1 _12825_ (.A1(_05501_),
    .A2(net563),
    .B1(_05827_),
    .B2(_05828_),
    .C1(_05751_),
    .X(_00760_));
 sky130_fd_sc_hd__xor2_1 _12826_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05789_),
    .X(_05829_));
 sky130_fd_sc_hd__and4_1 _12827_ (.A(_05807_),
    .B(_05821_),
    .C(_05817_),
    .D(_05826_),
    .X(_05830_));
 sky130_fd_sc_hd__o21a_1 _12828_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1(_05789_),
    .X(_05831_));
 sky130_fd_sc_hd__or4_1 _12829_ (.A(_05808_),
    .B(_05816_),
    .C(_05830_),
    .D(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__xor2_1 _12830_ (.A(_05829_),
    .B(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__mux2_1 _12831_ (.A0(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A1(_05833_),
    .S(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05834_));
 sky130_fd_sc_hd__and2_1 _12832_ (.A(_05652_),
    .B(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__clkbuf_1 _12833_ (.A(_05835_),
    .X(_00761_));
 sky130_fd_sc_hd__a22o_1 _12834_ (.A1(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_05789_),
    .B1(_05829_),
    .B2(_05832_),
    .X(_05836_));
 sky130_fd_sc_hd__xnor2_1 _12835_ (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05789_),
    .Y(_05837_));
 sky130_fd_sc_hd__xnor2_1 _12836_ (.A(_05836_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__or2_1 _12837_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05499_),
    .X(_05839_));
 sky130_fd_sc_hd__o211a_1 _12838_ (.A1(_05632_),
    .A2(_05838_),
    .B1(_05839_),
    .C1(_05675_),
    .X(_00762_));
 sky130_fd_sc_hd__and2_1 _12839_ (.A(_05490_),
    .B(_02310_),
    .X(_05840_));
 sky130_fd_sc_hd__clkbuf_1 _12840_ (.A(_05840_),
    .X(_00763_));
 sky130_fd_sc_hd__inv_2 _12841_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_05841_));
 sky130_fd_sc_hd__clkbuf_4 _12842_ (.A(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_4 _12843_ (.A(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__clkbuf_4 _12844_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05844_));
 sky130_fd_sc_hd__clkbuf_4 _12845_ (.A(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__or2_1 _12846_ (.A(net148),
    .B(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__o211a_1 _12847_ (.A1(_05843_),
    .A2(net281),
    .B1(_05495_),
    .C1(_05846_),
    .X(_00764_));
 sky130_fd_sc_hd__clkbuf_4 _12848_ (.A(_03619_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_2 _12849_ (.A(_05844_),
    .X(_05848_));
 sky130_fd_sc_hd__or2_1 _12850_ (.A(net140),
    .B(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__o211a_1 _12851_ (.A1(_05843_),
    .A2(net207),
    .B1(_05847_),
    .C1(_05849_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _12852_ (.A(net646),
    .B(_05848_),
    .X(_05850_));
 sky130_fd_sc_hd__o211a_1 _12853_ (.A1(_05843_),
    .A2(net204),
    .B1(_05847_),
    .C1(_05850_),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _12854_ (.A(net645),
    .B(_05848_),
    .X(_05851_));
 sky130_fd_sc_hd__o211a_1 _12855_ (.A1(_05843_),
    .A2(net167),
    .B1(_05847_),
    .C1(_05851_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _12856_ (.A(_05845_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(_05852_));
 sky130_fd_sc_hd__o211a_1 _12857_ (.A1(_05843_),
    .A2(net176),
    .B1(_05847_),
    .C1(_05852_),
    .X(_00768_));
 sky130_fd_sc_hd__buf_2 _12858_ (.A(_05844_),
    .X(_05853_));
 sky130_fd_sc_hd__clkbuf_4 _12859_ (.A(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__clkbuf_4 _12860_ (.A(_05844_),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _12861_ (.A(_05855_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .Y(_05856_));
 sky130_fd_sc_hd__o211a_1 _12862_ (.A1(_05854_),
    .A2(net435),
    .B1(_05847_),
    .C1(_05856_),
    .X(_00769_));
 sky130_fd_sc_hd__nand2_1 _12863_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .Y(_05857_));
 sky130_fd_sc_hd__or2_1 _12864_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(_05858_));
 sky130_fd_sc_hd__a21oi_1 _12865_ (.A1(_05857_),
    .A2(_05858_),
    .B1(_05567_),
    .Y(_05859_));
 sky130_fd_sc_hd__clkbuf_4 _12866_ (.A(_05841_),
    .X(_05860_));
 sky130_fd_sc_hd__a31o_1 _12867_ (.A1(_05567_),
    .A2(_05857_),
    .A3(_05858_),
    .B1(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__o221a_1 _12868_ (.A1(_05854_),
    .A2(net635),
    .B1(_05859_),
    .B2(_05861_),
    .C1(_05751_),
    .X(_00770_));
 sky130_fd_sc_hd__and3_1 _12869_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(_05862_));
 sky130_fd_sc_hd__a21oi_1 _12870_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .Y(_05863_));
 sky130_fd_sc_hd__or2_1 _12871_ (.A(_05862_),
    .B(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__nor2_1 _12872_ (.A(_05859_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21o_1 _12873_ (.A1(_05859_),
    .A2(_05864_),
    .B1(_05842_),
    .X(_05866_));
 sky130_fd_sc_hd__o221a_1 _12874_ (.A1(_05854_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B1(_05865_),
    .B2(_05866_),
    .C1(_05751_),
    .X(_00771_));
 sky130_fd_sc_hd__nand2_1 _12875_ (.A(_05566_),
    .B(_05862_),
    .Y(_05867_));
 sky130_fd_sc_hd__o31a_1 _12876_ (.A1(_05567_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A3(_05858_),
    .B1(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__and2_1 _12877_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__o21ai_1 _12878_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_05868_),
    .B1(_05845_),
    .Y(_05870_));
 sky130_fd_sc_hd__o221a_1 _12879_ (.A1(_05854_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B1(_05869_),
    .B2(_05870_),
    .C1(_05751_),
    .X(_00772_));
 sky130_fd_sc_hd__clkbuf_4 _12880_ (.A(_05853_),
    .X(_05871_));
 sky130_fd_sc_hd__or3_1 _12881_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .C(_05858_),
    .X(_05872_));
 sky130_fd_sc_hd__nand2_1 _12882_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_05862_),
    .Y(_05873_));
 sky130_fd_sc_hd__mux2_1 _12883_ (.A0(_05872_),
    .A1(_05873_),
    .S(_05566_),
    .X(_05874_));
 sky130_fd_sc_hd__and2_1 _12884_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__o21ai_1 _12885_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(_05874_),
    .B1(_05845_),
    .Y(_05876_));
 sky130_fd_sc_hd__o221a_1 _12886_ (.A1(_05871_),
    .A2(net553),
    .B1(_05875_),
    .B2(_05876_),
    .C1(_05751_),
    .X(_00773_));
 sky130_fd_sc_hd__inv_2 _12887_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_05877_));
 sky130_fd_sc_hd__clkbuf_4 _12888_ (.A(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__o21ai_1 _12889_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(_05872_),
    .B1(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__a31o_1 _12890_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A3(_05862_),
    .B1(_05878_),
    .X(_05880_));
 sky130_fd_sc_hd__inv_2 _12891_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .Y(_05881_));
 sky130_fd_sc_hd__a21oi_1 _12892_ (.A1(_05879_),
    .A2(_05880_),
    .B1(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__a31o_1 _12893_ (.A1(_05881_),
    .A2(_05879_),
    .A3(_05880_),
    .B1(_05860_),
    .X(_05883_));
 sky130_fd_sc_hd__o221a_1 _12894_ (.A1(_05871_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B1(_05882_),
    .B2(_05883_),
    .C1(_05751_),
    .X(_00774_));
 sky130_fd_sc_hd__and4_1 _12895_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .C(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .D(_05862_),
    .X(_05884_));
 sky130_fd_sc_hd__or3_1 _12896_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .C(_05872_),
    .X(_05885_));
 sky130_fd_sc_hd__inv_2 _12897_ (.A(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__mux2_1 _12898_ (.A0(_05884_),
    .A1(_05886_),
    .S(_05878_),
    .X(_05887_));
 sky130_fd_sc_hd__xnor2_1 _12899_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_1 _12900_ (.A(_05855_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__o211a_1 _12901_ (.A1(_05854_),
    .A2(net575),
    .B1(_05847_),
    .C1(_05889_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _12902_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_05885_),
    .X(_05890_));
 sky130_fd_sc_hd__nor2_1 _12903_ (.A(_05566_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__a31o_1 _12904_ (.A1(_05567_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A3(_05884_),
    .B1(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__xor2_1 _12905_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__or2_1 _12906_ (.A(_05848_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(_05894_));
 sky130_fd_sc_hd__o211a_1 _12907_ (.A1(_05843_),
    .A2(_05893_),
    .B1(_05894_),
    .C1(_05675_),
    .X(_00776_));
 sky130_fd_sc_hd__and3_1 _12908_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(_05884_),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_1 _12909_ (.A(_05566_),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__o31a_1 _12910_ (.A1(_05567_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A3(_05890_),
    .B1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__and2_1 _12911_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__o21ai_1 _12912_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_05897_),
    .B1(_05845_),
    .Y(_05899_));
 sky130_fd_sc_hd__o221a_1 _12913_ (.A1(_05871_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B1(_05898_),
    .B2(_05899_),
    .C1(_05751_),
    .X(_00777_));
 sky130_fd_sc_hd__nand3_1 _12914_ (.A(_05567_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_05895_),
    .Y(_05900_));
 sky130_fd_sc_hd__o41a_1 _12915_ (.A1(_05566_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A4(_05890_),
    .B1(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__nor2_1 _12916_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__a21o_1 _12917_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_05901_),
    .B1(_05842_),
    .X(_05903_));
 sky130_fd_sc_hd__o221a_1 _12918_ (.A1(_05871_),
    .A2(net557),
    .B1(_05902_),
    .B2(_05903_),
    .C1(_05751_),
    .X(_00778_));
 sky130_fd_sc_hd__or4_1 _12919_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .D(_05890_),
    .X(_05904_));
 sky130_fd_sc_hd__and3_1 _12920_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_05895_),
    .X(_05905_));
 sky130_fd_sc_hd__nand2_1 _12921_ (.A(_05567_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__o21a_1 _12922_ (.A1(_05567_),
    .A2(_05904_),
    .B1(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__and2_1 _12923_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__o21ai_1 _12924_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_05907_),
    .B1(_05845_),
    .Y(_05909_));
 sky130_fd_sc_hd__clkbuf_4 _12925_ (.A(_04538_),
    .X(_05910_));
 sky130_fd_sc_hd__o221a_1 _12926_ (.A1(_05871_),
    .A2(net627),
    .B1(_05908_),
    .B2(_05909_),
    .C1(_05910_),
    .X(_00779_));
 sky130_fd_sc_hd__nand3_1 _12927_ (.A(_05566_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_05905_),
    .Y(_05911_));
 sky130_fd_sc_hd__o31a_1 _12928_ (.A1(_05567_),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A3(_05904_),
    .B1(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__and2_1 _12929_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__o21ai_1 _12930_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_05912_),
    .B1(_05845_),
    .Y(_05914_));
 sky130_fd_sc_hd__o221a_1 _12931_ (.A1(_05871_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_05913_),
    .B2(_05914_),
    .C1(_05910_),
    .X(_00780_));
 sky130_fd_sc_hd__and3_1 _12932_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_05905_),
    .X(_05915_));
 sky130_fd_sc_hd__inv_2 _12933_ (.A(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__or3_1 _12934_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_05904_),
    .X(_05917_));
 sky130_fd_sc_hd__mux2_1 _12935_ (.A0(_05916_),
    .A1(_05917_),
    .S(_05878_),
    .X(_05918_));
 sky130_fd_sc_hd__nor2_1 _12936_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__a21o_1 _12937_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05918_),
    .B1(_05842_),
    .X(_05920_));
 sky130_fd_sc_hd__o221a_1 _12938_ (.A1(_05871_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_05919_),
    .B2(_05920_),
    .C1(_05910_),
    .X(_00781_));
 sky130_fd_sc_hd__o21a_1 _12939_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05917_),
    .B1(_05878_),
    .X(_05921_));
 sky130_fd_sc_hd__a21o_1 _12940_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_05915_),
    .B1(_05878_),
    .X(_05922_));
 sky130_fd_sc_hd__or2b_1 _12941_ (.A(_05921_),
    .B_N(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__nor2_1 _12942_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__a21o_1 _12943_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_05923_),
    .B1(_05842_),
    .X(_05925_));
 sky130_fd_sc_hd__o221a_1 _12944_ (.A1(_05871_),
    .A2(net467),
    .B1(_05924_),
    .B2(_05925_),
    .C1(_05910_),
    .X(_00782_));
 sky130_fd_sc_hd__a21oi_1 _12945_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_05922_),
    .B1(_05921_),
    .Y(_05926_));
 sky130_fd_sc_hd__clkbuf_4 _12946_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05927_));
 sky130_fd_sc_hd__buf_2 _12947_ (.A(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__or2_1 _12948_ (.A(_05848_),
    .B(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__o211a_1 _12949_ (.A1(_05843_),
    .A2(_05926_),
    .B1(_05929_),
    .C1(_05675_),
    .X(_00783_));
 sky130_fd_sc_hd__inv_2 _12950_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .Y(_05930_));
 sky130_fd_sc_hd__nor2_1 _12951_ (.A(_05930_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_05931_));
 sky130_fd_sc_hd__a21o_1 _12952_ (.A1(_05930_),
    .A2(net471),
    .B1(_05842_),
    .X(_05932_));
 sky130_fd_sc_hd__o221a_1 _12953_ (.A1(_05871_),
    .A2(net492),
    .B1(_05931_),
    .B2(_05932_),
    .C1(_05910_),
    .X(_00784_));
 sky130_fd_sc_hd__and2b_1 _12954_ (.A_N(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(_05933_));
 sky130_fd_sc_hd__xnor2_1 _12955_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__xnor2_1 _12956_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__xor2_1 _12957_ (.A(_05931_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__or2_1 _12958_ (.A(_05848_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_05937_));
 sky130_fd_sc_hd__clkbuf_4 _12959_ (.A(_04455_),
    .X(_05938_));
 sky130_fd_sc_hd__o211a_1 _12960_ (.A1(_05843_),
    .A2(_05936_),
    .B1(_05937_),
    .C1(_05938_),
    .X(_00785_));
 sky130_fd_sc_hd__and2_1 _12961_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_05934_),
    .X(_05939_));
 sky130_fd_sc_hd__nor2_1 _12962_ (.A(_05931_),
    .B(_05935_),
    .Y(_05940_));
 sky130_fd_sc_hd__o21ba_1 _12963_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1_N(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_05941_));
 sky130_fd_sc_hd__xnor2_1 _12964_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_05941_),
    .Y(_05942_));
 sky130_fd_sc_hd__or2_1 _12965_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__nand2_1 _12966_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_05942_),
    .Y(_05944_));
 sky130_fd_sc_hd__and2_1 _12967_ (.A(_05943_),
    .B(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__o21ai_2 _12968_ (.A1(_05939_),
    .A2(_05940_),
    .B1(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__o31a_1 _12969_ (.A1(_05939_),
    .A2(_05940_),
    .A3(_05945_),
    .B1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_05947_));
 sky130_fd_sc_hd__a22oi_1 _12970_ (.A1(_05860_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_05946_),
    .B2(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__and2b_1 _12971_ (.A_N(_05948_),
    .B(_03118_),
    .X(_05949_));
 sky130_fd_sc_hd__clkbuf_1 _12972_ (.A(_05949_),
    .X(_00786_));
 sky130_fd_sc_hd__o31a_1 _12973_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_05877_),
    .X(_05950_));
 sky130_fd_sc_hd__xnor2_1 _12974_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand2_1 _12975_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__or2_1 _12976_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_05951_),
    .X(_05953_));
 sky130_fd_sc_hd__and2_1 _12977_ (.A(_05952_),
    .B(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__nand2_1 _12978_ (.A(_05944_),
    .B(_05946_),
    .Y(_05955_));
 sky130_fd_sc_hd__xor2_1 _12979_ (.A(_05954_),
    .B(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__mux2_1 _12980_ (.A0(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_05956_),
    .S(_05844_),
    .X(_05957_));
 sky130_fd_sc_hd__and2_1 _12981_ (.A(_05652_),
    .B(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_1 _12982_ (.A(_05958_),
    .X(_00787_));
 sky130_fd_sc_hd__a21bo_1 _12983_ (.A1(_05944_),
    .A2(_05946_),
    .B1_N(_05954_),
    .X(_05959_));
 sky130_fd_sc_hd__nand2_1 _12984_ (.A(_05952_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__or4_1 _12985_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .C(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .D(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(_05961_));
 sky130_fd_sc_hd__nand2_1 _12986_ (.A(_05877_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__xor2_1 _12987_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__and2_1 _12988_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__nor2_1 _12989_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_05963_),
    .Y(_05965_));
 sky130_fd_sc_hd__or2_1 _12990_ (.A(_05964_),
    .B(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__xnor2_1 _12991_ (.A(_05960_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__or2_1 _12992_ (.A(_05848_),
    .B(net480),
    .X(_05968_));
 sky130_fd_sc_hd__o211a_1 _12993_ (.A1(_05843_),
    .A2(_05967_),
    .B1(_05968_),
    .C1(_05938_),
    .X(_00788_));
 sky130_fd_sc_hd__o21a_1 _12994_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(_05961_),
    .B1(_05877_),
    .X(_05969_));
 sky130_fd_sc_hd__xnor2_1 _12995_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__and2_1 _12996_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__or2_1 _12997_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_05970_),
    .X(_05972_));
 sky130_fd_sc_hd__or2b_1 _12998_ (.A(_05971_),
    .B_N(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__inv_2 _12999_ (.A(_05966_),
    .Y(_05974_));
 sky130_fd_sc_hd__a21o_1 _13000_ (.A1(_05960_),
    .A2(_05974_),
    .B1(_05964_),
    .X(_05975_));
 sky130_fd_sc_hd__and2_1 _13001_ (.A(_05973_),
    .B(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__o21ai_1 _13002_ (.A1(_05973_),
    .A2(_05975_),
    .B1(_05845_),
    .Y(_05977_));
 sky130_fd_sc_hd__o221a_1 _13003_ (.A1(_05871_),
    .A2(net411),
    .B1(_05976_),
    .B2(_05977_),
    .C1(_05910_),
    .X(_00789_));
 sky130_fd_sc_hd__inv_2 _13004_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .Y(_05978_));
 sky130_fd_sc_hd__or3_2 _13005_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .C(_05961_),
    .X(_05979_));
 sky130_fd_sc_hd__nor2_1 _13006_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05566_),
    .Y(_05980_));
 sky130_fd_sc_hd__nor2_1 _13007_ (.A(_05978_),
    .B(_05878_),
    .Y(_05981_));
 sky130_fd_sc_hd__a21oi_4 _13008_ (.A1(_05979_),
    .A2(_05980_),
    .B1(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_1 _13009_ (.A1(_05978_),
    .A2(_05979_),
    .B1(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__or2_1 _13010_ (.A(_05614_),
    .B(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__nand2_1 _13011_ (.A(_05614_),
    .B(_05983_),
    .Y(_05985_));
 sky130_fd_sc_hd__nand2_2 _13012_ (.A(_05984_),
    .B(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__a21oi_1 _13013_ (.A1(_05972_),
    .A2(_05975_),
    .B1(_05971_),
    .Y(_05987_));
 sky130_fd_sc_hd__nor2_1 _13014_ (.A(_05986_),
    .B(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__a21o_1 _13015_ (.A1(_05986_),
    .A2(_05987_),
    .B1(_05841_),
    .X(_05989_));
 sky130_fd_sc_hd__o2bb2a_1 _13016_ (.A1_N(_05841_),
    .A2_N(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_05988_),
    .B2(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__and2b_1 _13017_ (.A_N(_05990_),
    .B(_01512_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _13018_ (.A(_05991_),
    .X(_00790_));
 sky130_fd_sc_hd__nand2_1 _13019_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_05982_),
    .Y(_05992_));
 sky130_fd_sc_hd__or2_1 _13020_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_05982_),
    .X(_05993_));
 sky130_fd_sc_hd__nand2_1 _13021_ (.A(_05992_),
    .B(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__o21ai_1 _13022_ (.A1(_05986_),
    .A2(_05987_),
    .B1(_05984_),
    .Y(_05995_));
 sky130_fd_sc_hd__xnor2_1 _13023_ (.A(_05994_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__or2_1 _13024_ (.A(_05848_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(_05997_));
 sky130_fd_sc_hd__o211a_1 _13025_ (.A1(_05843_),
    .A2(_05996_),
    .B1(_05997_),
    .C1(_05938_),
    .X(_00791_));
 sky130_fd_sc_hd__clkbuf_4 _13026_ (.A(_05842_),
    .X(_05998_));
 sky130_fd_sc_hd__o21ai_1 _13027_ (.A1(_05964_),
    .A2(_05971_),
    .B1(_05972_),
    .Y(_05999_));
 sky130_fd_sc_hd__o311a_1 _13028_ (.A1(_05986_),
    .A2(_05999_),
    .A3(_05994_),
    .B1(_05992_),
    .C1(_05984_),
    .X(_06000_));
 sky130_fd_sc_hd__or2_1 _13029_ (.A(_05966_),
    .B(_05973_),
    .X(_06001_));
 sky130_fd_sc_hd__a2111o_1 _13030_ (.A1(_05952_),
    .A2(_05959_),
    .B1(_05986_),
    .C1(_06001_),
    .D1(_05994_),
    .X(_06002_));
 sky130_fd_sc_hd__buf_4 _13031_ (.A(_05982_),
    .X(_06003_));
 sky130_fd_sc_hd__xnor2_1 _13032_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__a21oi_2 _13033_ (.A1(_06000_),
    .A2(_06002_),
    .B1(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__and3_1 _13034_ (.A(_06004_),
    .B(_06000_),
    .C(_06002_),
    .X(_06006_));
 sky130_fd_sc_hd__nor2_1 _13035_ (.A(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__or2_1 _13036_ (.A(_05848_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_06008_));
 sky130_fd_sc_hd__o211a_1 _13037_ (.A1(_05998_),
    .A2(_06007_),
    .B1(_06008_),
    .C1(_05938_),
    .X(_00792_));
 sky130_fd_sc_hd__xnor2_1 _13038_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_05982_),
    .Y(_06009_));
 sky130_fd_sc_hd__clkbuf_4 _13039_ (.A(_06003_),
    .X(_06010_));
 sky130_fd_sc_hd__a21o_1 _13040_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_06010_),
    .B1(_06005_),
    .X(_06011_));
 sky130_fd_sc_hd__xnor2_1 _13041_ (.A(_06009_),
    .B(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__or2_1 _13042_ (.A(_05848_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_06013_));
 sky130_fd_sc_hd__o211a_1 _13043_ (.A1(_05998_),
    .A2(_06012_),
    .B1(_06013_),
    .C1(_05938_),
    .X(_00793_));
 sky130_fd_sc_hd__and2_1 _13044_ (.A(_05842_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(_06014_));
 sky130_fd_sc_hd__o21ai_1 _13045_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_06010_),
    .Y(_06015_));
 sky130_fd_sc_hd__o21ai_1 _13046_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_06010_),
    .B1(_06005_),
    .Y(_06016_));
 sky130_fd_sc_hd__xnor2_1 _13047_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_06003_),
    .Y(_06017_));
 sky130_fd_sc_hd__a21oi_1 _13048_ (.A1(_06015_),
    .A2(_06016_),
    .B1(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__a31o_1 _13049_ (.A1(_06017_),
    .A2(_06015_),
    .A3(_06016_),
    .B1(_05860_),
    .X(_06019_));
 sky130_fd_sc_hd__nor2_1 _13050_ (.A(_06018_),
    .B(_06019_),
    .Y(_06020_));
 sky130_fd_sc_hd__o21a_1 _13051_ (.A1(_06014_),
    .A2(_06020_),
    .B1(_04961_),
    .X(_00794_));
 sky130_fd_sc_hd__xnor2_1 _13052_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_06003_),
    .Y(_06021_));
 sky130_fd_sc_hd__a21o_1 _13053_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_06010_),
    .B1(_06018_),
    .X(_06022_));
 sky130_fd_sc_hd__xnor2_1 _13054_ (.A(_06021_),
    .B(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__or2_1 _13055_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_06024_));
 sky130_fd_sc_hd__o211a_1 _13056_ (.A1(_05998_),
    .A2(_06023_),
    .B1(_06024_),
    .C1(_05938_),
    .X(_00795_));
 sky130_fd_sc_hd__xnor2_1 _13057_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_06003_),
    .Y(_06025_));
 sky130_fd_sc_hd__nor3_1 _13058_ (.A(_06009_),
    .B(_06017_),
    .C(_06021_),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2_1 _13059_ (.A(_06005_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__o41ai_2 _13060_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A4(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_06003_),
    .Y(_06028_));
 sky130_fd_sc_hd__and2_1 _13061_ (.A(_06027_),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__xor2_1 _13062_ (.A(_06025_),
    .B(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__or2_1 _13063_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_06031_));
 sky130_fd_sc_hd__o211a_1 _13064_ (.A1(_05998_),
    .A2(_06030_),
    .B1(_06031_),
    .C1(_05938_),
    .X(_00796_));
 sky130_fd_sc_hd__xnor2_1 _13065_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_06003_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand2_1 _13066_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_06010_),
    .Y(_06033_));
 sky130_fd_sc_hd__o21ai_1 _13067_ (.A1(_06025_),
    .A2(_06029_),
    .B1(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__xnor2_1 _13068_ (.A(_06032_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__or2_1 _13069_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_06036_));
 sky130_fd_sc_hd__o211a_1 _13070_ (.A1(_05998_),
    .A2(_06035_),
    .B1(_06036_),
    .C1(_05938_),
    .X(_00797_));
 sky130_fd_sc_hd__xnor2_2 _13071_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06003_),
    .Y(_06037_));
 sky130_fd_sc_hd__or2_1 _13072_ (.A(_06025_),
    .B(_06032_),
    .X(_06038_));
 sky130_fd_sc_hd__o21ai_1 _13073_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_06003_),
    .Y(_06039_));
 sky130_fd_sc_hd__o21a_1 _13074_ (.A1(_06029_),
    .A2(_06038_),
    .B1(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__xor2_1 _13075_ (.A(_06037_),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__mux2_1 _13076_ (.A0(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A1(_06041_),
    .S(_05844_),
    .X(_06042_));
 sky130_fd_sc_hd__and2_1 _13077_ (.A(_05652_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__clkbuf_1 _13078_ (.A(_06043_),
    .X(_00798_));
 sky130_fd_sc_hd__xnor2_1 _13079_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_06003_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand2_1 _13080_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06010_),
    .Y(_06045_));
 sky130_fd_sc_hd__o21ai_1 _13081_ (.A1(_06037_),
    .A2(_06040_),
    .B1(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__xnor2_1 _13082_ (.A(_06044_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__or2_1 _13083_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(_06048_));
 sky130_fd_sc_hd__o211a_1 _13084_ (.A1(_05998_),
    .A2(_06047_),
    .B1(_06048_),
    .C1(_05938_),
    .X(_00799_));
 sky130_fd_sc_hd__and2_1 _13085_ (.A(_05842_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .X(_06049_));
 sky130_fd_sc_hd__or4_1 _13086_ (.A(_06027_),
    .B(_06037_),
    .C(_06038_),
    .D(_06044_),
    .X(_06050_));
 sky130_fd_sc_hd__o41ai_1 _13087_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A4(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_06010_),
    .Y(_06051_));
 sky130_fd_sc_hd__xnor2_1 _13088_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06010_),
    .Y(_06052_));
 sky130_fd_sc_hd__a31oi_2 _13089_ (.A1(_06028_),
    .A2(_06050_),
    .A3(net113),
    .B1(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__a41o_1 _13090_ (.A1(_06028_),
    .A2(_06052_),
    .A3(_06050_),
    .A4(net112),
    .B1(_05860_),
    .X(_06054_));
 sky130_fd_sc_hd__nor2_1 _13091_ (.A(_06053_),
    .B(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__o21a_1 _13092_ (.A1(_06049_),
    .A2(_06055_),
    .B1(_04961_),
    .X(_00800_));
 sky130_fd_sc_hd__a21o_1 _13093_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(_06010_),
    .B1(_06053_),
    .X(_06056_));
 sky130_fd_sc_hd__xnor2_1 _13094_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_06010_),
    .Y(_06057_));
 sky130_fd_sc_hd__xnor2_1 _13095_ (.A(_06056_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__or2_1 _13096_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06059_));
 sky130_fd_sc_hd__o211a_1 _13097_ (.A1(_05998_),
    .A2(_06058_),
    .B1(_06059_),
    .C1(_05938_),
    .X(_00801_));
 sky130_fd_sc_hd__and2_1 _13098_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_06060_));
 sky130_fd_sc_hd__nor2_1 _13099_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .Y(_06061_));
 sky130_fd_sc_hd__o21ai_1 _13100_ (.A1(_06060_),
    .A2(_06061_),
    .B1(_05855_),
    .Y(_06062_));
 sky130_fd_sc_hd__o211a_1 _13101_ (.A1(_05854_),
    .A2(net314),
    .B1(_05847_),
    .C1(_06062_),
    .X(_00802_));
 sky130_fd_sc_hd__and2b_1 _13102_ (.A_N(_05566_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_06063_));
 sky130_fd_sc_hd__xnor2_1 _13103_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xnor2_1 _13104_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nor2_1 _13105_ (.A(_06060_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__and2_1 _13106_ (.A(_06060_),
    .B(_06065_),
    .X(_06067_));
 sky130_fd_sc_hd__o21ai_1 _13107_ (.A1(_06066_),
    .A2(_06067_),
    .B1(_05855_),
    .Y(_06068_));
 sky130_fd_sc_hd__o211a_1 _13108_ (.A1(_05854_),
    .A2(net294),
    .B1(_05847_),
    .C1(_06068_),
    .X(_00803_));
 sky130_fd_sc_hd__clkbuf_4 _13109_ (.A(_01252_),
    .X(_06069_));
 sky130_fd_sc_hd__and2b_1 _13110_ (.A_N(_06064_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_06070_));
 sky130_fd_sc_hd__inv_2 _13111_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_06071_));
 sky130_fd_sc_hd__o21a_1 _13112_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_05877_),
    .X(_06072_));
 sky130_fd_sc_hd__xnor2_1 _13113_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__xnor2_1 _13114_ (.A(_06071_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__o21bai_2 _13115_ (.A1(_06070_),
    .A2(_06067_),
    .B1_N(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__or3b_1 _13116_ (.A(_06070_),
    .B(_06067_),
    .C_N(_06074_),
    .X(_06076_));
 sky130_fd_sc_hd__and2_1 _13117_ (.A(_05841_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .X(_06077_));
 sky130_fd_sc_hd__a31o_1 _13118_ (.A1(_05844_),
    .A2(_06075_),
    .A3(_06076_),
    .B1(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__and2_1 _13119_ (.A(_06069_),
    .B(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__clkbuf_1 _13120_ (.A(_06079_),
    .X(_00804_));
 sky130_fd_sc_hd__inv_2 _13121_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_06080_));
 sky130_fd_sc_hd__or2_1 _13122_ (.A(_06071_),
    .B(_06073_),
    .X(_06081_));
 sky130_fd_sc_hd__inv_2 _13123_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_06082_));
 sky130_fd_sc_hd__o31a_1 _13124_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B1(_05878_),
    .X(_06083_));
 sky130_fd_sc_hd__xnor2_1 _13125_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__nor2_1 _13126_ (.A(_06082_),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__and2_1 _13127_ (.A(_06082_),
    .B(_06084_),
    .X(_06086_));
 sky130_fd_sc_hd__or2_1 _13128_ (.A(_06085_),
    .B(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__and3_1 _13129_ (.A(_06081_),
    .B(_06075_),
    .C(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__a21oi_2 _13130_ (.A1(_06081_),
    .A2(_06075_),
    .B1(_06087_),
    .Y(_06089_));
 sky130_fd_sc_hd__or3_1 _13131_ (.A(_05841_),
    .B(_06088_),
    .C(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__o21a_1 _13132_ (.A1(_05844_),
    .A2(_06080_),
    .B1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__and2b_1 _13133_ (.A_N(_06091_),
    .B(_01512_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _13134_ (.A(_06092_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _13135_ (.A(_06085_),
    .B(_06089_),
    .X(_06093_));
 sky130_fd_sc_hd__or4_2 _13136_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .C(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .D(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_06094_));
 sky130_fd_sc_hd__nand2_1 _13137_ (.A(_05878_),
    .B(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__xor2_2 _13138_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__xnor2_2 _13139_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__xnor2_1 _13140_ (.A(_06093_),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _13141_ (.A(_05855_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__o211a_1 _13142_ (.A1(_05854_),
    .A2(net270),
    .B1(_05847_),
    .C1(_06099_),
    .X(_00806_));
 sky130_fd_sc_hd__inv_2 _13143_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .Y(_06100_));
 sky130_fd_sc_hd__o21a_1 _13144_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(_06094_),
    .B1(_05878_),
    .X(_06101_));
 sky130_fd_sc_hd__xnor2_1 _13145_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__nor2_2 _13146_ (.A(_06100_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__and2_1 _13147_ (.A(_06100_),
    .B(_06102_),
    .X(_06104_));
 sky130_fd_sc_hd__nor2_1 _13148_ (.A(_06103_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__and2b_1 _13149_ (.A_N(_06096_),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_06106_));
 sky130_fd_sc_hd__a21oi_1 _13150_ (.A1(_06093_),
    .A2(_06097_),
    .B1(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__xnor2_1 _13151_ (.A(_06105_),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__or2_1 _13152_ (.A(_05853_),
    .B(net539),
    .X(_06109_));
 sky130_fd_sc_hd__clkbuf_4 _13153_ (.A(_04455_),
    .X(_06110_));
 sky130_fd_sc_hd__o211a_1 _13154_ (.A1(_05998_),
    .A2(_06108_),
    .B1(_06109_),
    .C1(_06110_),
    .X(_00807_));
 sky130_fd_sc_hd__o31a_1 _13155_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A3(_06094_),
    .B1(_05877_),
    .X(_06111_));
 sky130_fd_sc_hd__mux2_2 _13156_ (.A0(_06111_),
    .A1(_05566_),
    .S(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06112_));
 sky130_fd_sc_hd__or4b_1 _13157_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(_06094_),
    .D_N(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06113_));
 sky130_fd_sc_hd__or2b_1 _13158_ (.A(_06112_),
    .B_N(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__and2_1 _13159_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__nor2_1 _13160_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_06114_),
    .Y(_06116_));
 sky130_fd_sc_hd__nor2_2 _13161_ (.A(_06115_),
    .B(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_1 _13162_ (.A(_06104_),
    .B(_06107_),
    .Y(_06118_));
 sky130_fd_sc_hd__nor2_1 _13163_ (.A(_06103_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__xnor2_1 _13164_ (.A(_06117_),
    .B(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_06120_),
    .S(_05844_),
    .X(_06121_));
 sky130_fd_sc_hd__and2_1 _13166_ (.A(_06069_),
    .B(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_1 _13167_ (.A(_06122_),
    .X(_00808_));
 sky130_fd_sc_hd__o21a_1 _13168_ (.A1(_06103_),
    .A2(_06118_),
    .B1(_06117_),
    .X(_06123_));
 sky130_fd_sc_hd__nand2_1 _13169_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_06112_),
    .Y(_06124_));
 sky130_fd_sc_hd__or2_1 _13170_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_06112_),
    .X(_06125_));
 sky130_fd_sc_hd__nand2_1 _13171_ (.A(_06124_),
    .B(_06125_),
    .Y(_06126_));
 sky130_fd_sc_hd__nor3_1 _13172_ (.A(_06115_),
    .B(_06123_),
    .C(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__o21ai_1 _13173_ (.A1(_06115_),
    .A2(_06123_),
    .B1(_06126_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_1 _13174_ (.A(_05845_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__o221a_1 _13175_ (.A1(_05855_),
    .A2(net388),
    .B1(_06127_),
    .B2(_06129_),
    .C1(_05910_),
    .X(_00809_));
 sky130_fd_sc_hd__o21ba_1 _13176_ (.A1(_06106_),
    .A2(_06103_),
    .B1_N(_06104_),
    .X(_06130_));
 sky130_fd_sc_hd__inv_2 _13177_ (.A(_06126_),
    .Y(_06131_));
 sky130_fd_sc_hd__or2b_1 _13178_ (.A(_06115_),
    .B_N(_06124_),
    .X(_06132_));
 sky130_fd_sc_hd__a32oi_4 _13179_ (.A1(_06117_),
    .A2(_06130_),
    .A3(_06131_),
    .B1(_06132_),
    .B2(_06125_),
    .Y(_06133_));
 sky130_fd_sc_hd__nor3b_1 _13180_ (.A(_06103_),
    .B(_06104_),
    .C_N(_06097_),
    .Y(_06134_));
 sky130_fd_sc_hd__o2111ai_4 _13181_ (.A1(_06085_),
    .A2(_06089_),
    .B1(_06117_),
    .C1(_06134_),
    .D1(_06131_),
    .Y(_06135_));
 sky130_fd_sc_hd__clkbuf_4 _13182_ (.A(_06112_),
    .X(_06136_));
 sky130_fd_sc_hd__xnor2_1 _13183_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__a21oi_2 _13184_ (.A1(_06133_),
    .A2(_06135_),
    .B1(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__and3_1 _13185_ (.A(_06137_),
    .B(_06133_),
    .C(_06135_),
    .X(_06139_));
 sky130_fd_sc_hd__o21ai_1 _13186_ (.A1(_06138_),
    .A2(_06139_),
    .B1(_05855_),
    .Y(_06140_));
 sky130_fd_sc_hd__o211a_1 _13187_ (.A1(_05854_),
    .A2(net494),
    .B1(_05847_),
    .C1(_06140_),
    .X(_00810_));
 sky130_fd_sc_hd__xor2_1 _13188_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_06136_),
    .X(_06141_));
 sky130_fd_sc_hd__clkbuf_4 _13189_ (.A(_06136_),
    .X(_06142_));
 sky130_fd_sc_hd__a21oi_1 _13190_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_06142_),
    .B1(_06138_),
    .Y(_06143_));
 sky130_fd_sc_hd__xnor2_1 _13191_ (.A(_06141_),
    .B(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__or2_1 _13192_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_06145_));
 sky130_fd_sc_hd__o211a_1 _13193_ (.A1(_05998_),
    .A2(_06144_),
    .B1(_06145_),
    .C1(_06110_),
    .X(_00811_));
 sky130_fd_sc_hd__o21a_1 _13194_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_06142_),
    .X(_06146_));
 sky130_fd_sc_hd__o21a_1 _13195_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_06142_),
    .B1(_06138_),
    .X(_06147_));
 sky130_fd_sc_hd__or2_1 _13196_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_06136_),
    .X(_06148_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_06136_),
    .Y(_06149_));
 sky130_fd_sc_hd__and2_1 _13198_ (.A(_06148_),
    .B(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__o21ai_2 _13199_ (.A1(_06146_),
    .A2(_06147_),
    .B1(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__o31a_1 _13200_ (.A1(_06150_),
    .A2(_06146_),
    .A3(_06147_),
    .B1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06152_));
 sky130_fd_sc_hd__a22o_1 _13201_ (.A1(_05860_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_06151_),
    .B2(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__and2_1 _13202_ (.A(_06069_),
    .B(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _13203_ (.A(_06154_),
    .X(_00812_));
 sky130_fd_sc_hd__xnor2_1 _13204_ (.A(_05930_),
    .B(_06136_),
    .Y(_06155_));
 sky130_fd_sc_hd__a21oi_1 _13205_ (.A1(_06149_),
    .A2(_06151_),
    .B1(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__a31o_1 _13206_ (.A1(_06149_),
    .A2(_06151_),
    .A3(_06155_),
    .B1(_05860_),
    .X(_06157_));
 sky130_fd_sc_hd__o221a_1 _13207_ (.A1(_05855_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_06156_),
    .B2(_06157_),
    .C1(_05910_),
    .X(_00813_));
 sky130_fd_sc_hd__nor2_1 _13208_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_06136_),
    .Y(_06158_));
 sky130_fd_sc_hd__nand2_1 _13209_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_06112_),
    .Y(_06159_));
 sky130_fd_sc_hd__and2b_1 _13210_ (.A_N(_06158_),
    .B(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__and4_1 _13211_ (.A(_06138_),
    .B(_06141_),
    .C(_06150_),
    .D(_06155_),
    .X(_06161_));
 sky130_fd_sc_hd__o41a_1 _13212_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A4(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_06142_),
    .X(_06162_));
 sky130_fd_sc_hd__or2_1 _13213_ (.A(_06161_),
    .B(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__or2_1 _13214_ (.A(_06160_),
    .B(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__nand2_1 _13215_ (.A(_06160_),
    .B(_06163_),
    .Y(_06165_));
 sky130_fd_sc_hd__and2_1 _13216_ (.A(_06164_),
    .B(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__or2_1 _13217_ (.A(_05853_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_06167_));
 sky130_fd_sc_hd__o211a_1 _13218_ (.A1(_05998_),
    .A2(_06166_),
    .B1(_06167_),
    .C1(_06110_),
    .X(_00814_));
 sky130_fd_sc_hd__xor2_1 _13219_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_06136_),
    .X(_06168_));
 sky130_fd_sc_hd__a21oi_1 _13220_ (.A1(_06159_),
    .A2(_06165_),
    .B1(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__a31o_1 _13221_ (.A1(_06159_),
    .A2(_06165_),
    .A3(_06168_),
    .B1(_05860_),
    .X(_06170_));
 sky130_fd_sc_hd__o221a_1 _13222_ (.A1(_05855_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_06169_),
    .B2(_06170_),
    .C1(_05910_),
    .X(_00815_));
 sky130_fd_sc_hd__nand2_1 _13223_ (.A(_05842_),
    .B(net489),
    .Y(_06171_));
 sky130_fd_sc_hd__o21a_1 _13224_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_06142_),
    .X(_06172_));
 sky130_fd_sc_hd__and2_1 _13225_ (.A(_06160_),
    .B(_06168_),
    .X(_06173_));
 sky130_fd_sc_hd__and2_1 _13226_ (.A(_06163_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__nor2_1 _13227_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06136_),
    .Y(_06175_));
 sky130_fd_sc_hd__nand2_1 _13228_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06136_),
    .Y(_06176_));
 sky130_fd_sc_hd__and2b_1 _13229_ (.A_N(_06175_),
    .B(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__o21ai_1 _13230_ (.A1(_06172_),
    .A2(_06174_),
    .B1(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__o31a_1 _13231_ (.A1(_06177_),
    .A2(_06172_),
    .A3(_06174_),
    .B1(_05844_),
    .X(_06179_));
 sky130_fd_sc_hd__nand2_1 _13232_ (.A(_06178_),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__a21boi_1 _13233_ (.A1(_06171_),
    .A2(_06180_),
    .B1_N(_01766_),
    .Y(_00816_));
 sky130_fd_sc_hd__xor2_1 _13234_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_06142_),
    .X(_06181_));
 sky130_fd_sc_hd__a21oi_1 _13235_ (.A1(_06176_),
    .A2(_06178_),
    .B1(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__a31o_1 _13236_ (.A1(_06176_),
    .A2(_06178_),
    .A3(_06181_),
    .B1(_05860_),
    .X(_06183_));
 sky130_fd_sc_hd__o221a_1 _13237_ (.A1(_05855_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_06182_),
    .B2(_06183_),
    .C1(_05910_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _13238_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06142_),
    .X(_06184_));
 sky130_fd_sc_hd__nand2_1 _13239_ (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06142_),
    .Y(_06185_));
 sky130_fd_sc_hd__nand2_1 _13240_ (.A(_06184_),
    .B(_06185_),
    .Y(_06186_));
 sky130_fd_sc_hd__and3_1 _13241_ (.A(_06177_),
    .B(_06173_),
    .C(_06181_),
    .X(_06187_));
 sky130_fd_sc_hd__o41a_1 _13242_ (.A1(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A3(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A4(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_06142_),
    .X(_06188_));
 sky130_fd_sc_hd__a211o_1 _13243_ (.A1(_06161_),
    .A2(_06187_),
    .B1(_06188_),
    .C1(_06162_),
    .X(_06189_));
 sky130_fd_sc_hd__xnor2_1 _13244_ (.A(_06186_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__mux2_1 _13245_ (.A0(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A1(_06190_),
    .S(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06191_));
 sky130_fd_sc_hd__and2_1 _13246_ (.A(_06069_),
    .B(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _13247_ (.A(_06192_),
    .X(_00818_));
 sky130_fd_sc_hd__or2b_1 _13248_ (.A(_06186_),
    .B_N(_06189_),
    .X(_06193_));
 sky130_fd_sc_hd__xnor2_1 _13249_ (.A(_05978_),
    .B(_06142_),
    .Y(_06194_));
 sky130_fd_sc_hd__a21oi_1 _13250_ (.A1(_06185_),
    .A2(_06193_),
    .B1(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__a31o_1 _13251_ (.A1(_06185_),
    .A2(_06193_),
    .A3(_06194_),
    .B1(_05860_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_4 _13252_ (.A(_04538_),
    .X(_06197_));
 sky130_fd_sc_hd__o221a_1 _13253_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_05854_),
    .B1(_06195_),
    .B2(_06196_),
    .C1(_06197_),
    .X(_00819_));
 sky130_fd_sc_hd__and2_1 _13254_ (.A(_05845_),
    .B(_01979_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_1 _13255_ (.A(_06198_),
    .X(_00820_));
 sky130_fd_sc_hd__inv_2 _13256_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_06199_));
 sky130_fd_sc_hd__clkbuf_4 _13257_ (.A(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_4 _13258_ (.A(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__clkbuf_4 _13259_ (.A(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_4 _13260_ (.A(_03619_),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_4 _13261_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06204_));
 sky130_fd_sc_hd__buf_2 _13262_ (.A(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__or2_1 _13263_ (.A(net647),
    .B(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__o211a_1 _13264_ (.A1(_06202_),
    .A2(net148),
    .B1(_06203_),
    .C1(_06206_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _13265_ (.A(net648),
    .B(_06205_),
    .X(_06207_));
 sky130_fd_sc_hd__o211a_1 _13266_ (.A1(_06202_),
    .A2(net140),
    .B1(_06203_),
    .C1(_06207_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _13267_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B(_06205_),
    .X(_06208_));
 sky130_fd_sc_hd__o211a_1 _13268_ (.A1(_06202_),
    .A2(net295),
    .B1(_06203_),
    .C1(_06208_),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _13269_ (.A(_06205_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(_06209_));
 sky130_fd_sc_hd__o211a_1 _13270_ (.A1(_06202_),
    .A2(net287),
    .B1(_06203_),
    .C1(_06209_),
    .X(_00824_));
 sky130_fd_sc_hd__clkbuf_4 _13271_ (.A(_06204_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_4 _13272_ (.A(_06204_),
    .X(_06211_));
 sky130_fd_sc_hd__nand2_1 _13273_ (.A(_06211_),
    .B(net456),
    .Y(_06212_));
 sky130_fd_sc_hd__o211a_1 _13274_ (.A1(_06210_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B1(_06203_),
    .C1(_06212_),
    .X(_00825_));
 sky130_fd_sc_hd__nand2_1 _13275_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .Y(_06213_));
 sky130_fd_sc_hd__or2_1 _13276_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(_06214_));
 sky130_fd_sc_hd__a21oi_1 _13277_ (.A1(_06213_),
    .A2(_06214_),
    .B1(_05928_),
    .Y(_06215_));
 sky130_fd_sc_hd__clkbuf_4 _13278_ (.A(_06200_),
    .X(_06216_));
 sky130_fd_sc_hd__a31o_1 _13279_ (.A1(_05928_),
    .A2(_06213_),
    .A3(_06214_),
    .B1(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__o221a_1 _13280_ (.A1(_06210_),
    .A2(net598),
    .B1(_06215_),
    .B2(_06217_),
    .C1(_06197_),
    .X(_00826_));
 sky130_fd_sc_hd__and3_1 _13281_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .C(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(_06218_));
 sky130_fd_sc_hd__a21oi_1 _13282_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .Y(_06219_));
 sky130_fd_sc_hd__or2_1 _13283_ (.A(_06218_),
    .B(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__nor2_1 _13284_ (.A(_06215_),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__a21o_1 _13285_ (.A1(_06215_),
    .A2(_06220_),
    .B1(_06201_),
    .X(_06222_));
 sky130_fd_sc_hd__o221a_1 _13286_ (.A1(_06210_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B1(_06221_),
    .B2(_06222_),
    .C1(_06197_),
    .X(_00827_));
 sky130_fd_sc_hd__clkbuf_4 _13287_ (.A(_06204_),
    .X(_06223_));
 sky130_fd_sc_hd__nand2_1 _13288_ (.A(_05928_),
    .B(_06218_),
    .Y(_06224_));
 sky130_fd_sc_hd__or3_1 _13289_ (.A(_05927_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(_06214_),
    .X(_06225_));
 sky130_fd_sc_hd__a21oi_1 _13290_ (.A1(_06224_),
    .A2(_06225_),
    .B1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .Y(_06226_));
 sky130_fd_sc_hd__a31o_1 _13291_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(_06224_),
    .A3(_06225_),
    .B1(_06216_),
    .X(_06227_));
 sky130_fd_sc_hd__o221a_1 _13292_ (.A1(_06223_),
    .A2(net516),
    .B1(_06226_),
    .B2(_06227_),
    .C1(_06197_),
    .X(_00828_));
 sky130_fd_sc_hd__or3_1 _13293_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(_06214_),
    .X(_06228_));
 sky130_fd_sc_hd__nand2_1 _13294_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_06218_),
    .Y(_06229_));
 sky130_fd_sc_hd__mux2_1 _13295_ (.A0(_06228_),
    .A1(_06229_),
    .S(_05927_),
    .X(_06230_));
 sky130_fd_sc_hd__and2_1 _13296_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__clkbuf_4 _13297_ (.A(_06204_),
    .X(_06232_));
 sky130_fd_sc_hd__o21ai_1 _13298_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_06230_),
    .B1(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__o221a_1 _13299_ (.A1(_06223_),
    .A2(net577),
    .B1(_06231_),
    .B2(_06233_),
    .C1(_06197_),
    .X(_00829_));
 sky130_fd_sc_hd__inv_2 _13300_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_06234_));
 sky130_fd_sc_hd__clkbuf_4 _13301_ (.A(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__o21ai_1 _13302_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(_06228_),
    .B1(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__a31o_1 _13303_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A3(_06218_),
    .B1(_06235_),
    .X(_06237_));
 sky130_fd_sc_hd__inv_2 _13304_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .Y(_06238_));
 sky130_fd_sc_hd__a21oi_1 _13305_ (.A1(_06236_),
    .A2(_06237_),
    .B1(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__a31o_1 _13306_ (.A1(_06238_),
    .A2(_06236_),
    .A3(_06237_),
    .B1(_06216_),
    .X(_06240_));
 sky130_fd_sc_hd__o221a_1 _13307_ (.A1(_06223_),
    .A2(net595),
    .B1(_06239_),
    .B2(_06240_),
    .C1(_06197_),
    .X(_00830_));
 sky130_fd_sc_hd__and4_1 _13308_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .C(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .D(_06218_),
    .X(_06241_));
 sky130_fd_sc_hd__or3_1 _13309_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .C(_06228_),
    .X(_06242_));
 sky130_fd_sc_hd__inv_2 _13310_ (.A(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__mux2_1 _13311_ (.A0(_06241_),
    .A1(_06243_),
    .S(_06235_),
    .X(_06244_));
 sky130_fd_sc_hd__xnor2_1 _13312_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_1 _13313_ (.A(_06232_),
    .B(_06245_),
    .Y(_06246_));
 sky130_fd_sc_hd__o211a_1 _13314_ (.A1(_06210_),
    .A2(net637),
    .B1(_06203_),
    .C1(_06246_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _13315_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_06242_),
    .X(_06247_));
 sky130_fd_sc_hd__nor2_1 _13316_ (.A(_05927_),
    .B(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__a31o_1 _13317_ (.A1(_05928_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A3(_06241_),
    .B1(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__xor2_1 _13318_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_2 _13319_ (.A(_06204_),
    .X(_06251_));
 sky130_fd_sc_hd__or2_1 _13320_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(_06252_));
 sky130_fd_sc_hd__o211a_1 _13321_ (.A1(_06202_),
    .A2(_06250_),
    .B1(_06252_),
    .C1(_06110_),
    .X(_00832_));
 sky130_fd_sc_hd__and3_1 _13322_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(_06241_),
    .X(_06253_));
 sky130_fd_sc_hd__nand2_1 _13323_ (.A(_05927_),
    .B(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__o31a_1 _13324_ (.A1(_05928_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A3(_06247_),
    .B1(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__and2_1 _13325_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__o21ai_1 _13326_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_06255_),
    .B1(_06232_),
    .Y(_06257_));
 sky130_fd_sc_hd__o221a_1 _13327_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_06256_),
    .B2(_06257_),
    .C1(_06197_),
    .X(_00833_));
 sky130_fd_sc_hd__nand3_1 _13328_ (.A(_05928_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_06253_),
    .Y(_06258_));
 sky130_fd_sc_hd__o41a_1 _13329_ (.A1(_05927_),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A3(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A4(_06247_),
    .B1(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__nor2_1 _13330_ (.A(net483),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__a21o_1 _13331_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A2(_06259_),
    .B1(_06201_),
    .X(_06261_));
 sky130_fd_sc_hd__o221a_1 _13332_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B1(_06260_),
    .B2(_06261_),
    .C1(_06197_),
    .X(_00834_));
 sky130_fd_sc_hd__or4_1 _13333_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .D(_06247_),
    .X(_06262_));
 sky130_fd_sc_hd__and3_1 _13334_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .C(_06253_),
    .X(_06263_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(_05928_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__o21a_1 _13336_ (.A1(_05928_),
    .A2(_06262_),
    .B1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__and2_1 _13337_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__o21ai_1 _13338_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_06265_),
    .B1(_06232_),
    .Y(_06267_));
 sky130_fd_sc_hd__o221a_1 _13339_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B1(_06266_),
    .B2(_06267_),
    .C1(_06197_),
    .X(_00835_));
 sky130_fd_sc_hd__inv_2 _13340_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .Y(_06268_));
 sky130_fd_sc_hd__and2_1 _13341_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_06263_),
    .X(_06269_));
 sky130_fd_sc_hd__nor2_1 _13342_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_06262_),
    .Y(_06270_));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(_06269_),
    .A1(_06270_),
    .S(_06235_),
    .X(_06271_));
 sky130_fd_sc_hd__a21oi_1 _13344_ (.A1(_06268_),
    .A2(_06271_),
    .B1(_06201_),
    .Y(_06272_));
 sky130_fd_sc_hd__o21ai_1 _13345_ (.A1(_06268_),
    .A2(_06271_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__o211a_1 _13346_ (.A1(_06210_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_06203_),
    .C1(_06273_),
    .X(_00836_));
 sky130_fd_sc_hd__nand2_1 _13347_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_06269_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand2_1 _13348_ (.A(_06268_),
    .B(_06270_),
    .Y(_06275_));
 sky130_fd_sc_hd__mux2_1 _13349_ (.A0(_06274_),
    .A1(_06275_),
    .S(_06235_),
    .X(_06276_));
 sky130_fd_sc_hd__nor2_1 _13350_ (.A(net568),
    .B(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__a21o_1 _13351_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_06276_),
    .B1(_06216_),
    .X(_06278_));
 sky130_fd_sc_hd__o221a_1 _13352_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B1(_06277_),
    .B2(_06278_),
    .C1(_06197_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _13353_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_06275_),
    .X(_06279_));
 sky130_fd_sc_hd__and3_1 _13354_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_06269_),
    .X(_06280_));
 sky130_fd_sc_hd__nand2_1 _13355_ (.A(_05927_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__o21a_1 _13356_ (.A1(_05928_),
    .A2(_06279_),
    .B1(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__and2_1 _13357_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__o21ai_1 _13358_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_06282_),
    .B1(_06232_),
    .Y(_06284_));
 sky130_fd_sc_hd__clkbuf_4 _13359_ (.A(_04538_),
    .X(_06285_));
 sky130_fd_sc_hd__o221a_1 _13360_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_06283_),
    .B2(_06284_),
    .C1(_06285_),
    .X(_00838_));
 sky130_fd_sc_hd__o21a_1 _13361_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_06279_),
    .B1(_06235_),
    .X(_06286_));
 sky130_fd_sc_hd__a21o_1 _13362_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_06280_),
    .B1(_06235_),
    .X(_06287_));
 sky130_fd_sc_hd__or2b_1 _13363_ (.A(_06286_),
    .B_N(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nor2_1 _13364_ (.A(net467),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__a21o_1 _13365_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_06288_),
    .B1(_06216_),
    .X(_06290_));
 sky130_fd_sc_hd__o221a_1 _13366_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B1(_06289_),
    .B2(_06290_),
    .C1(_06285_),
    .X(_00839_));
 sky130_fd_sc_hd__a21oi_1 _13367_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_06287_),
    .B1(_06286_),
    .Y(_06291_));
 sky130_fd_sc_hd__clkbuf_4 _13368_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_06292_));
 sky130_fd_sc_hd__clkbuf_4 _13369_ (.A(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__or2_1 _13370_ (.A(_06251_),
    .B(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__o211a_1 _13371_ (.A1(_06202_),
    .A2(_06291_),
    .B1(_06294_),
    .C1(_06110_),
    .X(_00840_));
 sky130_fd_sc_hd__inv_2 _13372_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .Y(_06295_));
 sky130_fd_sc_hd__nor2_1 _13373_ (.A(_06295_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_06296_));
 sky130_fd_sc_hd__a21o_1 _13374_ (.A1(_06295_),
    .A2(net610),
    .B1(_06216_),
    .X(_06297_));
 sky130_fd_sc_hd__o221a_1 _13375_ (.A1(_06223_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_06296_),
    .B2(net611),
    .C1(_06285_),
    .X(_00841_));
 sky130_fd_sc_hd__and2b_1 _13376_ (.A_N(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_06298_));
 sky130_fd_sc_hd__xnor2_1 _13377_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__xnor2_1 _13378_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__xor2_1 _13379_ (.A(_06296_),
    .B(_06300_),
    .X(_06301_));
 sky130_fd_sc_hd__or2_1 _13380_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_06302_));
 sky130_fd_sc_hd__o211a_1 _13381_ (.A1(_06202_),
    .A2(_06301_),
    .B1(_06302_),
    .C1(_06110_),
    .X(_00842_));
 sky130_fd_sc_hd__o21a_1 _13382_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_06235_),
    .X(_06303_));
 sky130_fd_sc_hd__xnor2_1 _13383_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__nor2_1 _13384_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__nand2_1 _13385_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_06304_),
    .Y(_06306_));
 sky130_fd_sc_hd__or2b_1 _13386_ (.A(_06305_),
    .B_N(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__nand2_1 _13387_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_06299_),
    .Y(_06308_));
 sky130_fd_sc_hd__o21a_1 _13388_ (.A1(_06296_),
    .A2(_06300_),
    .B1(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__a21o_1 _13389_ (.A1(_06307_),
    .A2(_06309_),
    .B1(_06199_),
    .X(_06310_));
 sky130_fd_sc_hd__nor2_1 _13390_ (.A(_06307_),
    .B(_06309_),
    .Y(_06311_));
 sky130_fd_sc_hd__a2bb2o_1 _13391_ (.A1_N(_06310_),
    .A2_N(_06311_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B2(_06200_),
    .X(_06312_));
 sky130_fd_sc_hd__and2_1 _13392_ (.A(_06069_),
    .B(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_1 _13393_ (.A(_06313_),
    .X(_00843_));
 sky130_fd_sc_hd__o31a_1 _13394_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A3(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_06235_),
    .X(_06314_));
 sky130_fd_sc_hd__xnor2_1 _13395_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__and2_1 _13396_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__or2_1 _13397_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_06315_),
    .X(_06317_));
 sky130_fd_sc_hd__and2b_1 _13398_ (.A_N(_06316_),
    .B(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__o21ai_1 _13399_ (.A1(_06305_),
    .A2(_06309_),
    .B1(_06306_),
    .Y(_06319_));
 sky130_fd_sc_hd__xor2_1 _13400_ (.A(_06318_),
    .B(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_06320_),
    .S(_06204_),
    .X(_06321_));
 sky130_fd_sc_hd__and2_1 _13402_ (.A(_06069_),
    .B(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__clkbuf_1 _13403_ (.A(_06322_),
    .X(_00844_));
 sky130_fd_sc_hd__a21o_1 _13404_ (.A1(_06317_),
    .A2(_06319_),
    .B1(_06316_),
    .X(_06323_));
 sky130_fd_sc_hd__or4_2 _13405_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .C(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .D(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_06324_));
 sky130_fd_sc_hd__nand2_1 _13406_ (.A(_06234_),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__xor2_1 _13407_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__and2_1 _13408_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__nor2_1 _13409_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_06326_),
    .Y(_06328_));
 sky130_fd_sc_hd__nor2_1 _13410_ (.A(_06327_),
    .B(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__xor2_1 _13411_ (.A(_06323_),
    .B(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__or2_1 _13412_ (.A(_06251_),
    .B(net512),
    .X(_06331_));
 sky130_fd_sc_hd__o211a_1 _13413_ (.A1(_06202_),
    .A2(_06330_),
    .B1(_06331_),
    .C1(_06110_),
    .X(_00845_));
 sky130_fd_sc_hd__nor2_1 _13414_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06324_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_1 _13415_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__or2_1 _13416_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_06334_));
 sky130_fd_sc_hd__nand2_1 _13417_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_05927_),
    .Y(_06335_));
 sky130_fd_sc_hd__o21a_1 _13418_ (.A1(_06332_),
    .A2(_06334_),
    .B1(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__buf_2 _13419_ (.A(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__nand3_2 _13420_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_06333_),
    .C(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__a21o_1 _13421_ (.A1(_06333_),
    .A2(_06337_),
    .B1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_06339_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(_06338_),
    .B(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__a21o_1 _13423_ (.A1(_06323_),
    .A2(_06329_),
    .B1(_06327_),
    .X(_06341_));
 sky130_fd_sc_hd__and2_1 _13424_ (.A(_06340_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__o21ai_1 _13425_ (.A1(_06340_),
    .A2(_06341_),
    .B1(_06205_),
    .Y(_06343_));
 sky130_fd_sc_hd__o221a_1 _13426_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B1(_06342_),
    .B2(_06343_),
    .C1(_06285_),
    .X(_00846_));
 sky130_fd_sc_hd__nand2_1 _13427_ (.A(_06339_),
    .B(_06341_),
    .Y(_06344_));
 sky130_fd_sc_hd__xnor2_1 _13428_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_06337_),
    .Y(_06345_));
 sky130_fd_sc_hd__a31o_1 _13429_ (.A1(_06338_),
    .A2(_06344_),
    .A3(_06345_),
    .B1(_06199_),
    .X(_06346_));
 sky130_fd_sc_hd__a21oi_1 _13430_ (.A1(_06338_),
    .A2(_06344_),
    .B1(_06345_),
    .Y(_06347_));
 sky130_fd_sc_hd__a2bb2o_1 _13431_ (.A1_N(_06346_),
    .A2_N(_06347_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B2(_06200_),
    .X(_06348_));
 sky130_fd_sc_hd__and2_1 _13432_ (.A(_06069_),
    .B(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__clkbuf_1 _13433_ (.A(_06349_),
    .X(_00847_));
 sky130_fd_sc_hd__xnor2_1 _13434_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_06337_),
    .Y(_06350_));
 sky130_fd_sc_hd__buf_4 _13435_ (.A(_06337_),
    .X(_06351_));
 sky130_fd_sc_hd__clkbuf_4 _13436_ (.A(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__a21o_1 _13437_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A2(_06352_),
    .B1(_06347_),
    .X(_06353_));
 sky130_fd_sc_hd__and2_1 _13438_ (.A(_06350_),
    .B(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__o21ai_1 _13439_ (.A1(_06350_),
    .A2(_06353_),
    .B1(_06205_),
    .Y(_06355_));
 sky130_fd_sc_hd__o221a_1 _13440_ (.A1(_06211_),
    .A2(net593),
    .B1(_06354_),
    .B2(_06355_),
    .C1(_06285_),
    .X(_00848_));
 sky130_fd_sc_hd__o21ai_1 _13441_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_06351_),
    .Y(_06356_));
 sky130_fd_sc_hd__and3_1 _13442_ (.A(_06329_),
    .B(_06338_),
    .C(_06339_),
    .X(_06357_));
 sky130_fd_sc_hd__nor2_1 _13443_ (.A(_06345_),
    .B(_06350_),
    .Y(_06358_));
 sky130_fd_sc_hd__or2b_1 _13444_ (.A(_06327_),
    .B_N(_06338_),
    .X(_06359_));
 sky130_fd_sc_hd__and3_1 _13445_ (.A(_06339_),
    .B(_06359_),
    .C(_06358_),
    .X(_06360_));
 sky130_fd_sc_hd__a31oi_2 _13446_ (.A1(_06323_),
    .A2(_06357_),
    .A3(_06358_),
    .B1(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__and2_1 _13447_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_06337_),
    .X(_06362_));
 sky130_fd_sc_hd__nor2_1 _13448_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_06337_),
    .Y(_06363_));
 sky130_fd_sc_hd__or2_1 _13449_ (.A(_06362_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__a21oi_2 _13450_ (.A1(_06356_),
    .A2(_06361_),
    .B1(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__and3_1 _13451_ (.A(_06364_),
    .B(_06356_),
    .C(_06361_),
    .X(_06366_));
 sky130_fd_sc_hd__nor2_1 _13452_ (.A(_06365_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__or2_1 _13453_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_06368_));
 sky130_fd_sc_hd__o211a_1 _13454_ (.A1(_06202_),
    .A2(_06367_),
    .B1(_06368_),
    .C1(_06110_),
    .X(_00849_));
 sky130_fd_sc_hd__xnor2_2 _13455_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_06351_),
    .Y(_06369_));
 sky130_fd_sc_hd__o21a_1 _13456_ (.A1(_06362_),
    .A2(_06365_),
    .B1(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__o31ai_1 _13457_ (.A1(_06362_),
    .A2(_06365_),
    .A3(_06369_),
    .B1(_06205_),
    .Y(_06371_));
 sky130_fd_sc_hd__o221a_1 _13458_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B1(_06370_),
    .B2(_06371_),
    .C1(_06285_),
    .X(_00850_));
 sky130_fd_sc_hd__nand2_1 _13459_ (.A(_06201_),
    .B(net409),
    .Y(_06372_));
 sky130_fd_sc_hd__o21a_1 _13460_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_06352_),
    .B1(_06365_),
    .X(_06373_));
 sky130_fd_sc_hd__o21a_1 _13461_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_06351_),
    .X(_06374_));
 sky130_fd_sc_hd__xnor2_1 _13462_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_06351_),
    .Y(_06375_));
 sky130_fd_sc_hd__o21ba_1 _13463_ (.A1(_06373_),
    .A2(_06374_),
    .B1_N(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__or3b_1 _13464_ (.A(_06374_),
    .B(_06373_),
    .C_N(_06375_),
    .X(_06377_));
 sky130_fd_sc_hd__or3b_1 _13465_ (.A(_06200_),
    .B(_06376_),
    .C_N(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__a21boi_1 _13466_ (.A1(_06372_),
    .A2(_06378_),
    .B1_N(_01766_),
    .Y(_00851_));
 sky130_fd_sc_hd__xnor2_1 _13467_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_06351_),
    .Y(_06379_));
 sky130_fd_sc_hd__a21o_1 _13468_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_06352_),
    .B1(_06376_),
    .X(_06380_));
 sky130_fd_sc_hd__xnor2_1 _13469_ (.A(_06379_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__or2_1 _13470_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_06382_));
 sky130_fd_sc_hd__o211a_1 _13471_ (.A1(_06202_),
    .A2(_06381_),
    .B1(_06382_),
    .C1(_06110_),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_1 _13472_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_06351_),
    .Y(_06383_));
 sky130_fd_sc_hd__nor3_1 _13473_ (.A(_06369_),
    .B(_06375_),
    .C(_06379_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_1 _13474_ (.A(_06365_),
    .B(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__o21a_1 _13475_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_06351_),
    .X(_06386_));
 sky130_fd_sc_hd__nor2_1 _13476_ (.A(_06374_),
    .B(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__and2_1 _13477_ (.A(_06385_),
    .B(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__nor2_1 _13478_ (.A(_06383_),
    .B(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__and2_1 _13479_ (.A(_06383_),
    .B(_06388_),
    .X(_06390_));
 sky130_fd_sc_hd__o21ai_1 _13480_ (.A1(_06389_),
    .A2(_06390_),
    .B1(_06232_),
    .Y(_06391_));
 sky130_fd_sc_hd__o211a_1 _13481_ (.A1(_06210_),
    .A2(net336),
    .B1(_06203_),
    .C1(_06391_),
    .X(_00853_));
 sky130_fd_sc_hd__a21o_1 _13482_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .A2(_06352_),
    .B1(_06389_),
    .X(_06392_));
 sky130_fd_sc_hd__xnor2_1 _13483_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_06337_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_1 _13484_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__a21o_1 _13485_ (.A1(_06392_),
    .A2(_06393_),
    .B1(_06216_),
    .X(_06395_));
 sky130_fd_sc_hd__o221a_1 _13486_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_06394_),
    .B2(_06395_),
    .C1(_06285_),
    .X(_00854_));
 sky130_fd_sc_hd__xnor2_1 _13487_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06351_),
    .Y(_06396_));
 sky130_fd_sc_hd__inv_2 _13488_ (.A(_06352_),
    .Y(_06397_));
 sky130_fd_sc_hd__nor2_1 _13489_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .Y(_06398_));
 sky130_fd_sc_hd__or2_1 _13490_ (.A(_06383_),
    .B(_06393_),
    .X(_06399_));
 sky130_fd_sc_hd__o22a_1 _13491_ (.A1(_06397_),
    .A2(_06398_),
    .B1(_06399_),
    .B2(_06388_),
    .X(_06400_));
 sky130_fd_sc_hd__xor2_1 _13492_ (.A(_06396_),
    .B(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__mux2_1 _13493_ (.A0(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A1(_06401_),
    .S(_06204_),
    .X(_06402_));
 sky130_fd_sc_hd__and2_1 _13494_ (.A(_06069_),
    .B(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _13495_ (.A(_06403_),
    .X(_00855_));
 sky130_fd_sc_hd__nand2_1 _13496_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06352_),
    .Y(_06404_));
 sky130_fd_sc_hd__o21ai_1 _13497_ (.A1(_06396_),
    .A2(_06400_),
    .B1(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__xnor2_2 _13498_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_06351_),
    .Y(_06406_));
 sky130_fd_sc_hd__nor2_1 _13499_ (.A(_06405_),
    .B(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__a21o_1 _13500_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06216_),
    .X(_06408_));
 sky130_fd_sc_hd__o221a_1 _13501_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B1(_06407_),
    .B2(_06408_),
    .C1(_06285_),
    .X(_00856_));
 sky130_fd_sc_hd__and2_1 _13502_ (.A(_06216_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .X(_06409_));
 sky130_fd_sc_hd__or4_1 _13503_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .C(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .D(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_06410_));
 sky130_fd_sc_hd__or3_1 _13504_ (.A(_06396_),
    .B(_06399_),
    .C(_06406_),
    .X(_06411_));
 sky130_fd_sc_hd__o2bb2a_1 _13505_ (.A1_N(_06352_),
    .A2_N(_06410_),
    .B1(_06411_),
    .B2(_06385_),
    .X(_06412_));
 sky130_fd_sc_hd__xnor2_1 _13506_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06352_),
    .Y(_06413_));
 sky130_fd_sc_hd__a21oi_1 _13507_ (.A1(_06387_),
    .A2(_06412_),
    .B1(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__a31o_1 _13508_ (.A1(_06387_),
    .A2(_06413_),
    .A3(_06412_),
    .B1(_06200_),
    .X(_06415_));
 sky130_fd_sc_hd__nor2_1 _13509_ (.A(_06414_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__o21a_1 _13510_ (.A1(_06409_),
    .A2(_06416_),
    .B1(_04961_),
    .X(_00857_));
 sky130_fd_sc_hd__a21o_1 _13511_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(_06352_),
    .B1(_06414_),
    .X(_06417_));
 sky130_fd_sc_hd__xnor2_1 _13512_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_06352_),
    .Y(_06418_));
 sky130_fd_sc_hd__xnor2_1 _13513_ (.A(_06417_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__or2_1 _13514_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06420_));
 sky130_fd_sc_hd__o211a_1 _13515_ (.A1(_06201_),
    .A2(_06419_),
    .B1(_06420_),
    .C1(_06110_),
    .X(_00858_));
 sky130_fd_sc_hd__and2_1 _13516_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_06421_));
 sky130_fd_sc_hd__nor2_1 _13517_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .Y(_06422_));
 sky130_fd_sc_hd__o21ai_1 _13518_ (.A1(_06421_),
    .A2(_06422_),
    .B1(_06232_),
    .Y(_06423_));
 sky130_fd_sc_hd__o211a_1 _13519_ (.A1(_06210_),
    .A2(net330),
    .B1(_06203_),
    .C1(_06423_),
    .X(_00859_));
 sky130_fd_sc_hd__and2b_1 _13520_ (.A_N(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_06424_));
 sky130_fd_sc_hd__xnor2_1 _13521_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__and2b_1 _13522_ (.A_N(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__and2b_1 _13523_ (.A_N(_06425_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_06427_));
 sky130_fd_sc_hd__nor2_1 _13524_ (.A(_06426_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__xnor2_1 _13525_ (.A(_06421_),
    .B(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__nand2_1 _13526_ (.A(_06232_),
    .B(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__o211a_1 _13527_ (.A1(_06210_),
    .A2(net299),
    .B1(_06203_),
    .C1(_06430_),
    .X(_00860_));
 sky130_fd_sc_hd__inv_2 _13528_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_06431_));
 sky130_fd_sc_hd__nor2_1 _13529_ (.A(_06232_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__nor2_1 _13530_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_06398_),
    .Y(_06433_));
 sky130_fd_sc_hd__xnor2_1 _13531_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__and2b_1 _13532_ (.A_N(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__and2b_1 _13533_ (.A_N(_06434_),
    .B(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .X(_06436_));
 sky130_fd_sc_hd__nor2_1 _13534_ (.A(_06435_),
    .B(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__a21o_1 _13535_ (.A1(_06421_),
    .A2(_06428_),
    .B1(_06427_),
    .X(_06438_));
 sky130_fd_sc_hd__o21ai_1 _13536_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06205_),
    .Y(_06439_));
 sky130_fd_sc_hd__a21oi_1 _13537_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__o21a_1 _13538_ (.A1(_06432_),
    .A2(_06440_),
    .B1(_04961_),
    .X(_00861_));
 sky130_fd_sc_hd__o31a_1 _13539_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A3(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_06235_),
    .X(_06441_));
 sky130_fd_sc_hd__xnor2_1 _13540_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__nor2_1 _13541_ (.A(_06080_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_06080_),
    .B(_06442_),
    .Y(_06444_));
 sky130_fd_sc_hd__or2b_1 _13543_ (.A(_06443_),
    .B_N(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__a21o_1 _13544_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06436_),
    .X(_06446_));
 sky130_fd_sc_hd__xnor2_1 _13545_ (.A(_06445_),
    .B(_06446_),
    .Y(_06447_));
 sky130_fd_sc_hd__mux2_1 _13546_ (.A0(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A1(_06447_),
    .S(_06204_),
    .X(_06448_));
 sky130_fd_sc_hd__and2_1 _13547_ (.A(_06069_),
    .B(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__clkbuf_1 _13548_ (.A(_06449_),
    .X(_00862_));
 sky130_fd_sc_hd__a21oi_2 _13549_ (.A1(_06444_),
    .A2(_06446_),
    .B1(_06443_),
    .Y(_06450_));
 sky130_fd_sc_hd__inv_2 _13550_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .Y(_06451_));
 sky130_fd_sc_hd__nand2_1 _13551_ (.A(_06234_),
    .B(_06410_),
    .Y(_06452_));
 sky130_fd_sc_hd__xor2_1 _13552_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__nor2_1 _13553_ (.A(_06451_),
    .B(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__and2_1 _13554_ (.A(_06451_),
    .B(_06453_),
    .X(_06455_));
 sky130_fd_sc_hd__or2_1 _13555_ (.A(_06454_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__xor2_1 _13556_ (.A(_06450_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__or2_1 _13557_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_06458_));
 sky130_fd_sc_hd__clkbuf_4 _13558_ (.A(_04455_),
    .X(_06459_));
 sky130_fd_sc_hd__o211a_1 _13559_ (.A1(_06201_),
    .A2(_06457_),
    .B1(_06458_),
    .C1(_06459_),
    .X(_00863_));
 sky130_fd_sc_hd__nor2_1 _13560_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06410_),
    .Y(_06460_));
 sky130_fd_sc_hd__and2_1 _13561_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__nor2_1 _13562_ (.A(_05927_),
    .B(_06460_),
    .Y(_06462_));
 sky130_fd_sc_hd__mux2_2 _13563_ (.A0(_06462_),
    .A1(_05927_),
    .S(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06463_));
 sky130_fd_sc_hd__o21a_1 _13564_ (.A1(_06461_),
    .A2(_06463_),
    .B1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_06464_));
 sky130_fd_sc_hd__or3_1 _13565_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_06461_),
    .C(_06463_),
    .X(_06465_));
 sky130_fd_sc_hd__or2b_1 _13566_ (.A(_06464_),
    .B_N(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__o21ba_1 _13567_ (.A1(_06450_),
    .A2(_06456_),
    .B1_N(_06454_),
    .X(_06467_));
 sky130_fd_sc_hd__xor2_1 _13568_ (.A(_06466_),
    .B(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__or2_1 _13569_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_06469_));
 sky130_fd_sc_hd__o211a_1 _13570_ (.A1(_06201_),
    .A2(_06468_),
    .B1(_06469_),
    .C1(_06459_),
    .X(_00864_));
 sky130_fd_sc_hd__or2_1 _13571_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_06463_),
    .X(_06470_));
 sky130_fd_sc_hd__nand2_1 _13572_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_06463_),
    .Y(_06471_));
 sky130_fd_sc_hd__nand2_1 _13573_ (.A(_06470_),
    .B(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__or2_1 _13574_ (.A(_06456_),
    .B(_06466_),
    .X(_06473_));
 sky130_fd_sc_hd__o21ai_1 _13575_ (.A1(_06454_),
    .A2(_06464_),
    .B1(_06465_),
    .Y(_06474_));
 sky130_fd_sc_hd__o21a_1 _13576_ (.A1(_06450_),
    .A2(_06473_),
    .B1(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__xor2_1 _13577_ (.A(_06472_),
    .B(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_06476_),
    .S(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06477_));
 sky130_fd_sc_hd__and2_1 _13579_ (.A(_06069_),
    .B(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__clkbuf_1 _13580_ (.A(_06478_),
    .X(_00865_));
 sky130_fd_sc_hd__or2_1 _13581_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_06463_),
    .X(_06479_));
 sky130_fd_sc_hd__nand2_1 _13582_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_06463_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand2_1 _13583_ (.A(_06479_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__o21a_1 _13584_ (.A1(_06472_),
    .A2(_06475_),
    .B1(_06471_),
    .X(_06482_));
 sky130_fd_sc_hd__xor2_1 _13585_ (.A(_06481_),
    .B(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__or2_1 _13586_ (.A(_06251_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_06484_));
 sky130_fd_sc_hd__o211a_1 _13587_ (.A1(_06201_),
    .A2(_06483_),
    .B1(_06484_),
    .C1(_06459_),
    .X(_00866_));
 sky130_fd_sc_hd__clkbuf_4 _13588_ (.A(_01765_),
    .X(_06485_));
 sky130_fd_sc_hd__o311a_1 _13589_ (.A1(_06472_),
    .A2(_06474_),
    .A3(_06481_),
    .B1(_06480_),
    .C1(_06471_),
    .X(_06486_));
 sky130_fd_sc_hd__or4_2 _13590_ (.A(_06450_),
    .B(_06472_),
    .C(_06473_),
    .D(_06481_),
    .X(_06487_));
 sky130_fd_sc_hd__buf_2 _13591_ (.A(_06463_),
    .X(_06488_));
 sky130_fd_sc_hd__or2_1 _13592_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__nand2_1 _13593_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_06488_),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_1 _13594_ (.A(_06489_),
    .B(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(_06486_),
    .A2(_06487_),
    .B1(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__and3_1 _13596_ (.A(_06491_),
    .B(_06486_),
    .C(_06487_),
    .X(_06493_));
 sky130_fd_sc_hd__o21ai_1 _13597_ (.A1(_06492_),
    .A2(_06493_),
    .B1(_06232_),
    .Y(_06494_));
 sky130_fd_sc_hd__o211a_1 _13598_ (.A1(_06210_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_06485_),
    .C1(_06494_),
    .X(_00867_));
 sky130_fd_sc_hd__a21o_1 _13599_ (.A1(_06486_),
    .A2(_06487_),
    .B1(_06491_),
    .X(_06495_));
 sky130_fd_sc_hd__nor2_1 _13600_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_06488_),
    .Y(_06496_));
 sky130_fd_sc_hd__nand2_1 _13601_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_06488_),
    .Y(_06497_));
 sky130_fd_sc_hd__and2b_1 _13602_ (.A_N(_06496_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__a21oi_1 _13603_ (.A1(_06490_),
    .A2(_06495_),
    .B1(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__a31o_1 _13604_ (.A1(_06490_),
    .A2(_06495_),
    .A3(_06498_),
    .B1(_06216_),
    .X(_06500_));
 sky130_fd_sc_hd__o221a_1 _13605_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B1(_06499_),
    .B2(_06500_),
    .C1(_06285_),
    .X(_00868_));
 sky130_fd_sc_hd__clkbuf_4 _13606_ (.A(_01252_),
    .X(_06501_));
 sky130_fd_sc_hd__or2_1 _13607_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_06488_),
    .X(_06502_));
 sky130_fd_sc_hd__nand2_1 _13608_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_06488_),
    .Y(_06503_));
 sky130_fd_sc_hd__and2_1 _13609_ (.A(_06502_),
    .B(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__o211a_1 _13610_ (.A1(_06495_),
    .A2(_06496_),
    .B1(_06497_),
    .C1(_06490_),
    .X(_06505_));
 sky130_fd_sc_hd__xnor2_1 _13611_ (.A(_06504_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__mux2_1 _13612_ (.A0(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A1(_06506_),
    .S(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06507_));
 sky130_fd_sc_hd__and2_1 _13613_ (.A(_06501_),
    .B(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__clkbuf_1 _13614_ (.A(_06508_),
    .X(_00869_));
 sky130_fd_sc_hd__or2b_1 _13615_ (.A(_06505_),
    .B_N(_06504_),
    .X(_06509_));
 sky130_fd_sc_hd__xor2_1 _13616_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_06488_),
    .X(_06510_));
 sky130_fd_sc_hd__a21oi_1 _13617_ (.A1(_06503_),
    .A2(_06509_),
    .B1(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__a31o_1 _13618_ (.A1(_06503_),
    .A2(_06509_),
    .A3(_06510_),
    .B1(_06200_),
    .X(_06512_));
 sky130_fd_sc_hd__o221a_1 _13619_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_06511_),
    .B2(_06512_),
    .C1(_06285_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _13620_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_06488_),
    .X(_06513_));
 sky130_fd_sc_hd__clkbuf_4 _13621_ (.A(_06488_),
    .X(_06514_));
 sky130_fd_sc_hd__nand2_1 _13622_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__and2_1 _13623_ (.A(_06513_),
    .B(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__and3_1 _13624_ (.A(_06498_),
    .B(_06504_),
    .C(_06510_),
    .X(_06517_));
 sky130_fd_sc_hd__o41ai_2 _13625_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A4(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_06514_),
    .Y(_06518_));
 sky130_fd_sc_hd__a21bo_1 _13626_ (.A1(_06492_),
    .A2(_06517_),
    .B1_N(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__xor2_1 _13627_ (.A(_06516_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__or2_1 _13628_ (.A(_06204_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_06521_));
 sky130_fd_sc_hd__o211a_1 _13629_ (.A1(_06201_),
    .A2(_06520_),
    .B1(_06521_),
    .C1(_06459_),
    .X(_00871_));
 sky130_fd_sc_hd__nand2_1 _13630_ (.A(_06516_),
    .B(_06519_),
    .Y(_06522_));
 sky130_fd_sc_hd__xor2_2 _13631_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_06514_),
    .X(_06523_));
 sky130_fd_sc_hd__a21oi_1 _13632_ (.A1(_06515_),
    .A2(_06522_),
    .B1(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__a31o_1 _13633_ (.A1(_06515_),
    .A2(_06522_),
    .A3(_06523_),
    .B1(_06200_),
    .X(_06525_));
 sky130_fd_sc_hd__clkbuf_4 _13634_ (.A(_01474_),
    .X(_06526_));
 sky130_fd_sc_hd__o221a_1 _13635_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_06524_),
    .B2(_06525_),
    .C1(_06526_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _13636_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06488_),
    .X(_06527_));
 sky130_fd_sc_hd__nand2_1 _13637_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06514_),
    .Y(_06528_));
 sky130_fd_sc_hd__and2_1 _13638_ (.A(_06527_),
    .B(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__o21a_1 _13639_ (.A1(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_06514_),
    .X(_06530_));
 sky130_fd_sc_hd__a31o_1 _13640_ (.A1(_06516_),
    .A2(_06519_),
    .A3(_06523_),
    .B1(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__xor2_1 _13641_ (.A(_06529_),
    .B(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__mux2_1 _13642_ (.A0(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A1(_06532_),
    .S(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06533_));
 sky130_fd_sc_hd__and2_1 _13643_ (.A(_06501_),
    .B(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__clkbuf_1 _13644_ (.A(_06534_),
    .X(_00873_));
 sky130_fd_sc_hd__a21boi_1 _13645_ (.A1(_06529_),
    .A2(_06531_),
    .B1_N(_06528_),
    .Y(_06535_));
 sky130_fd_sc_hd__xor2_1 _13646_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_06514_),
    .X(_06536_));
 sky130_fd_sc_hd__and2_1 _13647_ (.A(_06535_),
    .B(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__o21ai_1 _13648_ (.A1(_06535_),
    .A2(_06536_),
    .B1(_06205_),
    .Y(_06538_));
 sky130_fd_sc_hd__o221a_1 _13649_ (.A1(_06211_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B1(_06537_),
    .B2(_06538_),
    .C1(_06526_),
    .X(_00874_));
 sky130_fd_sc_hd__and4_1 _13650_ (.A(_06516_),
    .B(_06523_),
    .C(_06529_),
    .D(_06536_),
    .X(_06539_));
 sky130_fd_sc_hd__nand3_1 _13651_ (.A(_06492_),
    .B(_06517_),
    .C(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2_1 _13652_ (.A(_06324_),
    .B(_06514_),
    .Y(_06541_));
 sky130_fd_sc_hd__or2_1 _13653_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06514_),
    .X(_06542_));
 sky130_fd_sc_hd__nand2_1 _13654_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06514_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand2_1 _13655_ (.A(_06542_),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__a31o_1 _13656_ (.A1(_06518_),
    .A2(_06540_),
    .A3(_06541_),
    .B1(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__a41oi_1 _13657_ (.A1(_06518_),
    .A2(_06544_),
    .A3(_06540_),
    .A4(_06541_),
    .B1(_06199_),
    .Y(_06546_));
 sky130_fd_sc_hd__a22o_1 _13658_ (.A1(_06200_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B1(_06545_),
    .B2(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__and2_1 _13659_ (.A(_06501_),
    .B(_06547_),
    .X(_06548_));
 sky130_fd_sc_hd__clkbuf_1 _13660_ (.A(_06548_),
    .X(_00875_));
 sky130_fd_sc_hd__xor2_1 _13661_ (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_06514_),
    .X(_06549_));
 sky130_fd_sc_hd__a21oi_1 _13662_ (.A1(_06543_),
    .A2(_06545_),
    .B1(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__a31o_1 _13663_ (.A1(_06543_),
    .A2(_06545_),
    .A3(_06549_),
    .B1(_06200_),
    .X(_06551_));
 sky130_fd_sc_hd__o221a_1 _13664_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_06210_),
    .B1(_06550_),
    .B2(_06551_),
    .C1(_06526_),
    .X(_00876_));
 sky130_fd_sc_hd__and2_1 _13665_ (.A(_06205_),
    .B(_01979_),
    .X(_06552_));
 sky130_fd_sc_hd__clkbuf_1 _13666_ (.A(_06552_),
    .X(_00877_));
 sky130_fd_sc_hd__buf_4 _13667_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06553_));
 sky130_fd_sc_hd__inv_2 _13668_ (.A(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__clkbuf_4 _13669_ (.A(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__buf_2 _13670_ (.A(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__buf_2 _13671_ (.A(_06553_),
    .X(_06557_));
 sky130_fd_sc_hd__or2_1 _13672_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__o211a_1 _13673_ (.A1(_06556_),
    .A2(net212),
    .B1(_06485_),
    .C1(_06558_),
    .X(_00878_));
 sky130_fd_sc_hd__or2_1 _13674_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .B(_06557_),
    .X(_06559_));
 sky130_fd_sc_hd__o211a_1 _13675_ (.A1(_06556_),
    .A2(net220),
    .B1(_06485_),
    .C1(_06559_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _13676_ (.A(_06557_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_06560_));
 sky130_fd_sc_hd__o211a_1 _13677_ (.A1(_06556_),
    .A2(net288),
    .B1(_06485_),
    .C1(_06560_),
    .X(_00880_));
 sky130_fd_sc_hd__clkbuf_4 _13678_ (.A(_06557_),
    .X(_06561_));
 sky130_fd_sc_hd__clkbuf_4 _13679_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .X(_06562_));
 sky130_fd_sc_hd__clkbuf_4 _13680_ (.A(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__nand2_1 _13681_ (.A(_06563_),
    .B(net453),
    .Y(_06564_));
 sky130_fd_sc_hd__o211a_1 _13682_ (.A1(_06561_),
    .A2(net403),
    .B1(_06485_),
    .C1(_06564_),
    .X(_00881_));
 sky130_fd_sc_hd__clkbuf_4 _13683_ (.A(_06562_),
    .X(_06565_));
 sky130_fd_sc_hd__nand2_1 _13684_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .Y(_06566_));
 sky130_fd_sc_hd__or2_1 _13685_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(_06567_));
 sky130_fd_sc_hd__a21oi_1 _13686_ (.A1(_06566_),
    .A2(_06567_),
    .B1(_06293_),
    .Y(_06568_));
 sky130_fd_sc_hd__clkbuf_4 _13687_ (.A(_06554_),
    .X(_06569_));
 sky130_fd_sc_hd__a31o_1 _13688_ (.A1(_06293_),
    .A2(_06566_),
    .A3(_06567_),
    .B1(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__o221a_1 _13689_ (.A1(_06565_),
    .A2(net524),
    .B1(_06568_),
    .B2(_06570_),
    .C1(_06526_),
    .X(_00882_));
 sky130_fd_sc_hd__and3_1 _13690_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .C(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(_06571_));
 sky130_fd_sc_hd__a21oi_1 _13691_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .Y(_06572_));
 sky130_fd_sc_hd__or2_1 _13692_ (.A(_06571_),
    .B(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__nor2_1 _13693_ (.A(_06568_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__a21o_1 _13694_ (.A1(_06568_),
    .A2(_06573_),
    .B1(_06555_),
    .X(_06575_));
 sky130_fd_sc_hd__o221a_1 _13695_ (.A1(_06565_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B1(_06574_),
    .B2(_06575_),
    .C1(_06526_),
    .X(_00883_));
 sky130_fd_sc_hd__nand2_1 _13696_ (.A(_06293_),
    .B(_06571_),
    .Y(_06576_));
 sky130_fd_sc_hd__or3_1 _13697_ (.A(_06292_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .C(_06567_),
    .X(_06577_));
 sky130_fd_sc_hd__a21oi_1 _13698_ (.A1(_06576_),
    .A2(_06577_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .Y(_06578_));
 sky130_fd_sc_hd__a31o_1 _13699_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_06576_),
    .A3(_06577_),
    .B1(_06569_),
    .X(_06579_));
 sky130_fd_sc_hd__o221a_1 _13700_ (.A1(_06565_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B1(_06578_),
    .B2(_06579_),
    .C1(_06526_),
    .X(_00884_));
 sky130_fd_sc_hd__or3_1 _13701_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .C(_06567_),
    .X(_06580_));
 sky130_fd_sc_hd__nand2_1 _13702_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_06571_),
    .Y(_06581_));
 sky130_fd_sc_hd__mux2_1 _13703_ (.A0(_06580_),
    .A1(_06581_),
    .S(_06292_),
    .X(_06582_));
 sky130_fd_sc_hd__and2_1 _13704_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(_06582_),
    .X(_06583_));
 sky130_fd_sc_hd__clkbuf_4 _13705_ (.A(_06562_),
    .X(_06584_));
 sky130_fd_sc_hd__o21ai_1 _13706_ (.A1(net516),
    .A2(_06582_),
    .B1(_06584_),
    .Y(_06585_));
 sky130_fd_sc_hd__o221a_1 _13707_ (.A1(_06565_),
    .A2(net590),
    .B1(_06583_),
    .B2(_06585_),
    .C1(_06526_),
    .X(_00885_));
 sky130_fd_sc_hd__inv_2 _13708_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .Y(_06586_));
 sky130_fd_sc_hd__clkbuf_4 _13709_ (.A(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__o21ai_1 _13710_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(_06580_),
    .B1(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__a31o_1 _13711_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A3(_06571_),
    .B1(_06587_),
    .X(_06589_));
 sky130_fd_sc_hd__inv_2 _13712_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .Y(_06590_));
 sky130_fd_sc_hd__a21oi_1 _13713_ (.A1(_06588_),
    .A2(_06589_),
    .B1(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__a31o_1 _13714_ (.A1(_06590_),
    .A2(_06588_),
    .A3(_06589_),
    .B1(_06569_),
    .X(_06592_));
 sky130_fd_sc_hd__o221a_1 _13715_ (.A1(_06565_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B1(_06591_),
    .B2(_06592_),
    .C1(_06526_),
    .X(_00886_));
 sky130_fd_sc_hd__and4_1 _13716_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .C(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .D(_06571_),
    .X(_06593_));
 sky130_fd_sc_hd__or3_1 _13717_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .C(_06580_),
    .X(_06594_));
 sky130_fd_sc_hd__inv_2 _13718_ (.A(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__mux2_1 _13719_ (.A0(_06593_),
    .A1(_06595_),
    .S(_06587_),
    .X(_06596_));
 sky130_fd_sc_hd__xnor2_1 _13720_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_06596_),
    .Y(_06597_));
 sky130_fd_sc_hd__nand2_1 _13721_ (.A(_06563_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__o211a_1 _13722_ (.A1(_06561_),
    .A2(net490),
    .B1(_06485_),
    .C1(_06598_),
    .X(_00887_));
 sky130_fd_sc_hd__or2_1 _13723_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_06594_),
    .X(_06599_));
 sky130_fd_sc_hd__and2_1 _13724_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_06593_),
    .X(_06600_));
 sky130_fd_sc_hd__nand2_1 _13725_ (.A(_06292_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__o21a_1 _13726_ (.A1(_06293_),
    .A2(_06599_),
    .B1(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__o21ai_1 _13727_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_06602_),
    .B1(_06562_),
    .Y(_06603_));
 sky130_fd_sc_hd__a21o_1 _13728_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_06602_),
    .B1(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__o211a_1 _13729_ (.A1(_06561_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B1(_06485_),
    .C1(_06604_),
    .X(_00888_));
 sky130_fd_sc_hd__nor2_1 _13730_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_06599_),
    .Y(_06605_));
 sky130_fd_sc_hd__nor2_1 _13731_ (.A(_06293_),
    .B(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__a21oi_2 _13732_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_06600_),
    .B1(_06587_),
    .Y(_06607_));
 sky130_fd_sc_hd__o21a_1 _13733_ (.A1(_06606_),
    .A2(_06607_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(_06608_));
 sky130_fd_sc_hd__o31ai_1 _13734_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_06606_),
    .A3(_06607_),
    .B1(_06584_),
    .Y(_06609_));
 sky130_fd_sc_hd__o221a_1 _13735_ (.A1(_06565_),
    .A2(net576),
    .B1(_06608_),
    .B2(_06609_),
    .C1(_06526_),
    .X(_00889_));
 sky130_fd_sc_hd__inv_2 _13736_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .Y(_06610_));
 sky130_fd_sc_hd__nand2_1 _13737_ (.A(_06610_),
    .B(_06605_),
    .Y(_06611_));
 sky130_fd_sc_hd__mux2_1 _13738_ (.A0(_06610_),
    .A1(_06611_),
    .S(_06587_),
    .X(_06612_));
 sky130_fd_sc_hd__o21a_1 _13739_ (.A1(_06607_),
    .A2(_06612_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(_06613_));
 sky130_fd_sc_hd__o31ai_1 _13740_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_06607_),
    .A3(_06612_),
    .B1(_06584_),
    .Y(_06614_));
 sky130_fd_sc_hd__o221a_1 _13741_ (.A1(_06565_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B1(_06613_),
    .B2(_06614_),
    .C1(_06526_),
    .X(_00890_));
 sky130_fd_sc_hd__and4_1 _13742_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .C(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .D(_06600_),
    .X(_06615_));
 sky130_fd_sc_hd__or2_1 _13743_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_06611_),
    .X(_06616_));
 sky130_fd_sc_hd__inv_2 _13744_ (.A(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__mux2_1 _13745_ (.A0(_06615_),
    .A1(_06617_),
    .S(_06587_),
    .X(_06618_));
 sky130_fd_sc_hd__xnor2_1 _13746_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__nand2_1 _13747_ (.A(_06563_),
    .B(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__o211a_1 _13748_ (.A1(_06561_),
    .A2(net597),
    .B1(_06485_),
    .C1(_06620_),
    .X(_00891_));
 sky130_fd_sc_hd__nand3_1 _13749_ (.A(_06292_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_06615_),
    .Y(_06621_));
 sky130_fd_sc_hd__o31a_1 _13750_ (.A1(_06292_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .A3(_06616_),
    .B1(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__o21ai_1 _13751_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_06622_),
    .B1(_06562_),
    .Y(_06623_));
 sky130_fd_sc_hd__a21o_1 _13752_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_06622_),
    .B1(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__o211a_1 _13753_ (.A1(_06561_),
    .A2(net561),
    .B1(_06485_),
    .C1(_06624_),
    .X(_00892_));
 sky130_fd_sc_hd__and3_1 _13754_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_06615_),
    .X(_06625_));
 sky130_fd_sc_hd__inv_2 _13755_ (.A(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__or3_1 _13756_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_06616_),
    .X(_06627_));
 sky130_fd_sc_hd__mux2_1 _13757_ (.A0(_06626_),
    .A1(_06627_),
    .S(_06587_),
    .X(_06628_));
 sky130_fd_sc_hd__nor2_1 _13758_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__a21o_1 _13759_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_06628_),
    .B1(_06569_),
    .X(_06630_));
 sky130_fd_sc_hd__clkbuf_4 _13760_ (.A(_01474_),
    .X(_06631_));
 sky130_fd_sc_hd__o221a_1 _13761_ (.A1(_06565_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B1(_06629_),
    .B2(_06630_),
    .C1(_06631_),
    .X(_00893_));
 sky130_fd_sc_hd__or2_1 _13762_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_06627_),
    .X(_06632_));
 sky130_fd_sc_hd__nor2_1 _13763_ (.A(_06293_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__a31o_1 _13764_ (.A1(_06293_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A3(_06625_),
    .B1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__xor2_1 _13765_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__or2_1 _13766_ (.A(_06557_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(_06636_));
 sky130_fd_sc_hd__o211a_1 _13767_ (.A1(_06556_),
    .A2(_06635_),
    .B1(_06636_),
    .C1(_06459_),
    .X(_00894_));
 sky130_fd_sc_hd__and3_1 _13768_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .C(_06625_),
    .X(_06637_));
 sky130_fd_sc_hd__nand2_1 _13769_ (.A(_06293_),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__o31a_1 _13770_ (.A1(_06293_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_06632_),
    .B1(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__and2_1 _13771_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__o21ai_1 _13772_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_06639_),
    .B1(_06584_),
    .Y(_06641_));
 sky130_fd_sc_hd__o221a_1 _13773_ (.A1(_06565_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .B1(_06640_),
    .B2(_06641_),
    .C1(_06631_),
    .X(_00895_));
 sky130_fd_sc_hd__o31a_1 _13774_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_06632_),
    .B1(_06587_),
    .X(_06642_));
 sky130_fd_sc_hd__a21oi_1 _13775_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_06637_),
    .B1(_06587_),
    .Y(_06643_));
 sky130_fd_sc_hd__o21a_1 _13776_ (.A1(_06642_),
    .A2(_06643_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_06644_));
 sky130_fd_sc_hd__o31ai_1 _13777_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_06642_),
    .A3(_06643_),
    .B1(_06584_),
    .Y(_06645_));
 sky130_fd_sc_hd__o221a_1 _13778_ (.A1(_06563_),
    .A2(net442),
    .B1(_06644_),
    .B2(_06645_),
    .C1(_06631_),
    .X(_00896_));
 sky130_fd_sc_hd__clkbuf_4 _13779_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_06646_));
 sky130_fd_sc_hd__clkbuf_4 _13780_ (.A(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__and2b_1 _13781_ (.A_N(_06643_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(_06648_));
 sky130_fd_sc_hd__o21ai_2 _13782_ (.A1(_06642_),
    .A2(_06648_),
    .B1(_06584_),
    .Y(_06649_));
 sky130_fd_sc_hd__o211a_1 _13783_ (.A1(_06561_),
    .A2(_06647_),
    .B1(_06485_),
    .C1(_06649_),
    .X(_00897_));
 sky130_fd_sc_hd__inv_2 _13784_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .Y(_06650_));
 sky130_fd_sc_hd__nor2_1 _13785_ (.A(_06650_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_06651_));
 sky130_fd_sc_hd__a21o_1 _13786_ (.A1(_06650_),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_06569_),
    .X(_06652_));
 sky130_fd_sc_hd__o221a_1 _13787_ (.A1(_06563_),
    .A2(net600),
    .B1(_06651_),
    .B2(_06652_),
    .C1(_06631_),
    .X(_00898_));
 sky130_fd_sc_hd__and2b_1 _13788_ (.A_N(_06292_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(_06653_));
 sky130_fd_sc_hd__xnor2_1 _13789_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__xnor2_1 _13790_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__xor2_1 _13791_ (.A(_06651_),
    .B(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__or2_1 _13792_ (.A(_06557_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_06657_));
 sky130_fd_sc_hd__o211a_1 _13793_ (.A1(_06556_),
    .A2(_06656_),
    .B1(_06657_),
    .C1(_06459_),
    .X(_00899_));
 sky130_fd_sc_hd__and2_1 _13794_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_06654_),
    .X(_06658_));
 sky130_fd_sc_hd__nor2_1 _13795_ (.A(_06651_),
    .B(_06655_),
    .Y(_06659_));
 sky130_fd_sc_hd__o21ba_1 _13796_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1_N(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_06660_));
 sky130_fd_sc_hd__xnor2_1 _13797_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__or2_1 _13798_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__nand2_1 _13799_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_06661_),
    .Y(_06663_));
 sky130_fd_sc_hd__and2_1 _13800_ (.A(_06662_),
    .B(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__o21ai_2 _13801_ (.A1(_06658_),
    .A2(_06659_),
    .B1(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__o31a_1 _13802_ (.A1(_06658_),
    .A2(_06659_),
    .A3(_06664_),
    .B1(_06553_),
    .X(_06666_));
 sky130_fd_sc_hd__a22oi_1 _13803_ (.A1(_06554_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_06665_),
    .B2(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__and2b_1 _13804_ (.A_N(_06667_),
    .B(_01512_),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_1 _13805_ (.A(_06668_),
    .X(_00900_));
 sky130_fd_sc_hd__o31a_1 _13806_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A3(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_06586_),
    .X(_06669_));
 sky130_fd_sc_hd__xnor2_1 _13807_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__or2_1 _13809_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_06670_),
    .X(_06672_));
 sky130_fd_sc_hd__and2_1 _13810_ (.A(_06671_),
    .B(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__nand2_1 _13811_ (.A(_06663_),
    .B(_06665_),
    .Y(_06674_));
 sky130_fd_sc_hd__xor2_1 _13812_ (.A(_06673_),
    .B(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__mux2_1 _13813_ (.A0(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .A1(_06675_),
    .S(_06562_),
    .X(_06676_));
 sky130_fd_sc_hd__and2_1 _13814_ (.A(_06501_),
    .B(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__clkbuf_1 _13815_ (.A(_06677_),
    .X(_00901_));
 sky130_fd_sc_hd__buf_4 _13816_ (.A(_01765_),
    .X(_06678_));
 sky130_fd_sc_hd__a21bo_1 _13817_ (.A1(_06663_),
    .A2(_06665_),
    .B1_N(_06673_),
    .X(_06679_));
 sky130_fd_sc_hd__nor4_1 _13818_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .C(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .D(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .Y(_06680_));
 sky130_fd_sc_hd__nand2_1 _13819_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__or2_1 _13820_ (.A(_06292_),
    .B(_06680_),
    .X(_06682_));
 sky130_fd_sc_hd__mux2_1 _13821_ (.A0(_06682_),
    .A1(_06586_),
    .S(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_06683_));
 sky130_fd_sc_hd__clkbuf_4 _13822_ (.A(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__and3_1 _13823_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_06681_),
    .C(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__a21oi_1 _13824_ (.A1(_06681_),
    .A2(_06684_),
    .B1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .Y(_06686_));
 sky130_fd_sc_hd__or2_1 _13825_ (.A(_06685_),
    .B(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__a21oi_2 _13826_ (.A1(_06671_),
    .A2(_06679_),
    .B1(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__and3_1 _13827_ (.A(_06671_),
    .B(_06679_),
    .C(_06687_),
    .X(_06689_));
 sky130_fd_sc_hd__o21ai_1 _13828_ (.A1(_06688_),
    .A2(_06689_),
    .B1(_06584_),
    .Y(_06690_));
 sky130_fd_sc_hd__o211a_1 _13829_ (.A1(_06561_),
    .A2(net639),
    .B1(_06678_),
    .C1(_06690_),
    .X(_00902_));
 sky130_fd_sc_hd__xnor2_2 _13830_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_06684_),
    .Y(_06691_));
 sky130_fd_sc_hd__o21a_1 _13831_ (.A1(_06685_),
    .A2(_06688_),
    .B1(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__o31ai_1 _13832_ (.A1(_06685_),
    .A2(_06688_),
    .A3(_06691_),
    .B1(_06584_),
    .Y(_06693_));
 sky130_fd_sc_hd__o221a_1 _13833_ (.A1(_06563_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B1(_06692_),
    .B2(_06693_),
    .C1(_06631_),
    .X(_00903_));
 sky130_fd_sc_hd__and2_1 _13834_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_06684_),
    .X(_06694_));
 sky130_fd_sc_hd__nor2_1 _13835_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_06684_),
    .Y(_06695_));
 sky130_fd_sc_hd__nor2_1 _13836_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__inv_2 _13837_ (.A(_06691_),
    .Y(_06697_));
 sky130_fd_sc_hd__a21o_1 _13838_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(_06684_),
    .B1(_06685_),
    .X(_06698_));
 sky130_fd_sc_hd__a21oi_1 _13839_ (.A1(_06688_),
    .A2(_06697_),
    .B1(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__xnor2_1 _13840_ (.A(_06696_),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__mux2_1 _13841_ (.A0(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A1(_06700_),
    .S(_06562_),
    .X(_06701_));
 sky130_fd_sc_hd__and2_1 _13842_ (.A(_06501_),
    .B(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_1 _13843_ (.A(_06702_),
    .X(_00904_));
 sky130_fd_sc_hd__xor2_1 _13844_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_06684_),
    .X(_06703_));
 sky130_fd_sc_hd__o21bai_1 _13845_ (.A1(_06695_),
    .A2(_06699_),
    .B1_N(_06694_),
    .Y(_06704_));
 sky130_fd_sc_hd__xnor2_1 _13846_ (.A(_06703_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_1 _13847_ (.A(_06563_),
    .B(_06705_),
    .Y(_06706_));
 sky130_fd_sc_hd__o211a_1 _13848_ (.A1(_06561_),
    .A2(net599),
    .B1(_06678_),
    .C1(_06706_),
    .X(_00905_));
 sky130_fd_sc_hd__buf_4 _13849_ (.A(_06684_),
    .X(_06707_));
 sky130_fd_sc_hd__xor2_1 _13850_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__nand2_1 _13851_ (.A(_06696_),
    .B(_06703_),
    .Y(_06709_));
 sky130_fd_sc_hd__a2111o_1 _13852_ (.A1(_06671_),
    .A2(_06679_),
    .B1(_06687_),
    .C1(_06691_),
    .D1(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a211oi_1 _13853_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(_06707_),
    .B1(_06694_),
    .C1(_06698_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_1 _13854_ (.A(_06710_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__xor2_1 _13855_ (.A(_06708_),
    .B(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__or2_1 _13856_ (.A(_06557_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(_06714_));
 sky130_fd_sc_hd__o211a_1 _13857_ (.A1(_06556_),
    .A2(_06713_),
    .B1(_06714_),
    .C1(_06459_),
    .X(_00906_));
 sky130_fd_sc_hd__xnor2_1 _13858_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_06707_),
    .Y(_06715_));
 sky130_fd_sc_hd__buf_2 _13859_ (.A(_06707_),
    .X(_06716_));
 sky130_fd_sc_hd__a21bo_1 _13860_ (.A1(_06710_),
    .A2(_06711_),
    .B1_N(_06708_),
    .X(_06717_));
 sky130_fd_sc_hd__a21bo_1 _13861_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_06716_),
    .B1_N(_06717_),
    .X(_06718_));
 sky130_fd_sc_hd__xnor2_1 _13862_ (.A(_06715_),
    .B(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__or2_1 _13863_ (.A(_06557_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_06720_));
 sky130_fd_sc_hd__o211a_1 _13864_ (.A1(_06556_),
    .A2(_06719_),
    .B1(_06720_),
    .C1(_06459_),
    .X(_00907_));
 sky130_fd_sc_hd__o21a_1 _13865_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_06707_),
    .X(_06721_));
 sky130_fd_sc_hd__o21ba_1 _13866_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_06716_),
    .B1_N(_06717_),
    .X(_06722_));
 sky130_fd_sc_hd__xnor2_1 _13867_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_06707_),
    .Y(_06723_));
 sky130_fd_sc_hd__or3b_1 _13868_ (.A(_06721_),
    .B(_06722_),
    .C_N(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__nand2_1 _13869_ (.A(_06553_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__o21ba_1 _13870_ (.A1(_06722_),
    .A2(_06721_),
    .B1_N(_06723_),
    .X(_06726_));
 sky130_fd_sc_hd__a2bb2o_1 _13871_ (.A1_N(_06725_),
    .A2_N(_06726_),
    .B1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B2(_06554_),
    .X(_06727_));
 sky130_fd_sc_hd__and2_1 _13872_ (.A(_06501_),
    .B(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_1 _13873_ (.A(_06728_),
    .X(_00908_));
 sky130_fd_sc_hd__xnor2_1 _13874_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_06707_),
    .Y(_06729_));
 sky130_fd_sc_hd__a21o_1 _13875_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_06716_),
    .B1(_06726_),
    .X(_06730_));
 sky130_fd_sc_hd__xnor2_1 _13876_ (.A(_06729_),
    .B(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__buf_2 _13877_ (.A(_06562_),
    .X(_06732_));
 sky130_fd_sc_hd__or2_1 _13878_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_06733_));
 sky130_fd_sc_hd__o211a_1 _13879_ (.A1(_06556_),
    .A2(_06731_),
    .B1(_06733_),
    .C1(_06459_),
    .X(_00909_));
 sky130_fd_sc_hd__nand2_1 _13880_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_06684_),
    .Y(_06734_));
 sky130_fd_sc_hd__or2_1 _13881_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_06684_),
    .X(_06735_));
 sky130_fd_sc_hd__nand2_1 _13882_ (.A(_06734_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__or3_1 _13883_ (.A(_06715_),
    .B(_06723_),
    .C(_06729_),
    .X(_06737_));
 sky130_fd_sc_hd__o21a_1 _13884_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_06716_),
    .X(_06738_));
 sky130_fd_sc_hd__nor2_1 _13885_ (.A(_06721_),
    .B(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__o21a_1 _13886_ (.A1(_06717_),
    .A2(_06737_),
    .B1(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__xor2_1 _13887_ (.A(_06736_),
    .B(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__or2_1 _13888_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_06742_));
 sky130_fd_sc_hd__o211a_1 _13889_ (.A1(_06556_),
    .A2(_06741_),
    .B1(_06742_),
    .C1(_06459_),
    .X(_00910_));
 sky130_fd_sc_hd__xnor2_2 _13890_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_06707_),
    .Y(_06743_));
 sky130_fd_sc_hd__o21ai_1 _13891_ (.A1(_06736_),
    .A2(_06740_),
    .B1(_06734_),
    .Y(_06744_));
 sky130_fd_sc_hd__xnor2_1 _13892_ (.A(_06743_),
    .B(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__or2_1 _13893_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_06746_));
 sky130_fd_sc_hd__clkbuf_4 _13894_ (.A(_04455_),
    .X(_06747_));
 sky130_fd_sc_hd__o211a_1 _13895_ (.A1(_06556_),
    .A2(_06745_),
    .B1(_06746_),
    .C1(_06747_),
    .X(_00911_));
 sky130_fd_sc_hd__xor2_1 _13896_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06707_),
    .X(_06748_));
 sky130_fd_sc_hd__o21a_1 _13897_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_06716_),
    .X(_06749_));
 sky130_fd_sc_hd__nor3_1 _13898_ (.A(_06736_),
    .B(_06740_),
    .C(_06743_),
    .Y(_06750_));
 sky130_fd_sc_hd__o31ai_1 _13899_ (.A1(_06748_),
    .A2(_06749_),
    .A3(_06750_),
    .B1(_06553_),
    .Y(_06751_));
 sky130_fd_sc_hd__o21a_1 _13900_ (.A1(_06749_),
    .A2(_06750_),
    .B1(_06748_),
    .X(_06752_));
 sky130_fd_sc_hd__a2bb2o_1 _13901_ (.A1_N(_06751_),
    .A2_N(_06752_),
    .B1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B2(_06554_),
    .X(_06753_));
 sky130_fd_sc_hd__and2_1 _13902_ (.A(_06501_),
    .B(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_1 _13903_ (.A(_06754_),
    .X(_00912_));
 sky130_fd_sc_hd__xnor2_1 _13904_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_06707_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21o_1 _13905_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_06716_),
    .B1(_06752_),
    .X(_06756_));
 sky130_fd_sc_hd__xnor2_1 _13906_ (.A(_06755_),
    .B(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__or2_1 _13907_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(_06758_));
 sky130_fd_sc_hd__o211a_1 _13908_ (.A1(_06555_),
    .A2(_06757_),
    .B1(_06758_),
    .C1(_06747_),
    .X(_00913_));
 sky130_fd_sc_hd__or2_1 _13909_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06716_),
    .X(_06759_));
 sky130_fd_sc_hd__nand2_1 _13910_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06716_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(_06759_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__or3b_1 _13912_ (.A(_06736_),
    .B(_06743_),
    .C_N(_06748_),
    .X(_06762_));
 sky130_fd_sc_hd__or4_1 _13913_ (.A(_06717_),
    .B(_06737_),
    .C(_06755_),
    .D(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__o21a_1 _13914_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_06716_),
    .X(_06764_));
 sky130_fd_sc_hd__nor2_1 _13915_ (.A(_06749_),
    .B(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__and3_1 _13916_ (.A(_06739_),
    .B(_06763_),
    .C(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__xor2_1 _13917_ (.A(_06761_),
    .B(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__mux2_1 _13918_ (.A0(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A1(_06767_),
    .S(_06553_),
    .X(_06768_));
 sky130_fd_sc_hd__and2_1 _13919_ (.A(_06501_),
    .B(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__clkbuf_1 _13920_ (.A(_06769_),
    .X(_00914_));
 sky130_fd_sc_hd__o21ai_1 _13921_ (.A1(_06761_),
    .A2(_06766_),
    .B1(_06760_),
    .Y(_06770_));
 sky130_fd_sc_hd__xnor2_1 _13922_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_06716_),
    .Y(_06771_));
 sky130_fd_sc_hd__xnor2_1 _13923_ (.A(_06770_),
    .B(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__or2_1 _13924_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06773_));
 sky130_fd_sc_hd__o211a_1 _13925_ (.A1(_06555_),
    .A2(_06772_),
    .B1(_06773_),
    .C1(_06747_),
    .X(_00915_));
 sky130_fd_sc_hd__and2_1 _13926_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_06774_));
 sky130_fd_sc_hd__nor2_1 _13927_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .Y(_06775_));
 sky130_fd_sc_hd__o21ai_1 _13928_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06584_),
    .Y(_06776_));
 sky130_fd_sc_hd__o211a_1 _13929_ (.A1(_06561_),
    .A2(net324),
    .B1(_06678_),
    .C1(_06776_),
    .X(_00916_));
 sky130_fd_sc_hd__and2b_1 _13930_ (.A_N(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_06777_));
 sky130_fd_sc_hd__xnor2_1 _13931_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__and2b_1 _13932_ (.A_N(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__and2b_1 _13933_ (.A_N(_06778_),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_06780_));
 sky130_fd_sc_hd__nor2_1 _13934_ (.A(_06779_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__xor2_1 _13935_ (.A(_06774_),
    .B(_06781_),
    .X(_06782_));
 sky130_fd_sc_hd__or2_1 _13936_ (.A(_06732_),
    .B(net578),
    .X(_06783_));
 sky130_fd_sc_hd__o211a_1 _13937_ (.A1(_06555_),
    .A2(_06782_),
    .B1(_06783_),
    .C1(_06747_),
    .X(_00917_));
 sky130_fd_sc_hd__o21a_1 _13938_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_06586_),
    .X(_06784_));
 sky130_fd_sc_hd__xnor2_1 _13939_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__and2_1 _13940_ (.A(_06431_),
    .B(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__nor2_1 _13941_ (.A(_06431_),
    .B(_06785_),
    .Y(_06787_));
 sky130_fd_sc_hd__nor2_1 _13942_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__a21o_1 _13943_ (.A1(_06774_),
    .A2(_06781_),
    .B1(_06780_),
    .X(_06789_));
 sky130_fd_sc_hd__nand2_1 _13944_ (.A(_06788_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__o21a_1 _13945_ (.A1(_06788_),
    .A2(_06789_),
    .B1(_06553_),
    .X(_06791_));
 sky130_fd_sc_hd__a22o_1 _13946_ (.A1(_06554_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .B1(_06790_),
    .B2(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__and2_1 _13947_ (.A(_06501_),
    .B(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__clkbuf_1 _13948_ (.A(_06793_),
    .X(_00918_));
 sky130_fd_sc_hd__inv_2 _13949_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_06794_));
 sky130_fd_sc_hd__o31a_1 _13950_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A3(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B1(_06587_),
    .X(_06795_));
 sky130_fd_sc_hd__xnor2_1 _13951_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__nor2_1 _13952_ (.A(_06794_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__nand2_1 _13953_ (.A(_06794_),
    .B(_06796_),
    .Y(_06798_));
 sky130_fd_sc_hd__or2b_1 _13954_ (.A(_06797_),
    .B_N(_06798_),
    .X(_06799_));
 sky130_fd_sc_hd__a21o_1 _13955_ (.A1(_06788_),
    .A2(_06789_),
    .B1(_06787_),
    .X(_06800_));
 sky130_fd_sc_hd__xnor2_1 _13956_ (.A(_06799_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__mux2_1 _13957_ (.A0(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .A1(_06801_),
    .S(_06553_),
    .X(_06802_));
 sky130_fd_sc_hd__and2_1 _13958_ (.A(_06501_),
    .B(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__clkbuf_1 _13959_ (.A(_06803_),
    .X(_00919_));
 sky130_fd_sc_hd__a21o_1 _13960_ (.A1(_06798_),
    .A2(_06800_),
    .B1(_06797_),
    .X(_06804_));
 sky130_fd_sc_hd__nor4_1 _13961_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .D(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .Y(_06805_));
 sky130_fd_sc_hd__nor2_1 _13962_ (.A(_06292_),
    .B(net116),
    .Y(_06806_));
 sky130_fd_sc_hd__mux2_2 _13963_ (.A0(_06806_),
    .A1(_06292_),
    .S(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_06807_));
 sky130_fd_sc_hd__a21o_1 _13964_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A2(net116),
    .B1(_06807_),
    .X(_06808_));
 sky130_fd_sc_hd__and2_1 _13965_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_06808_),
    .X(_06809_));
 sky130_fd_sc_hd__or2_1 _13966_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_06808_),
    .X(_06810_));
 sky130_fd_sc_hd__nor2b_1 _13967_ (.A(_06809_),
    .B_N(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__xor2_1 _13968_ (.A(_06804_),
    .B(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__or2_1 _13969_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_06813_));
 sky130_fd_sc_hd__o211a_1 _13970_ (.A1(_06555_),
    .A2(_06812_),
    .B1(_06813_),
    .C1(_06747_),
    .X(_00920_));
 sky130_fd_sc_hd__and2_1 _13971_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_06807_),
    .X(_06814_));
 sky130_fd_sc_hd__or2_1 _13972_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_06807_),
    .X(_06815_));
 sky130_fd_sc_hd__and2b_1 _13973_ (.A_N(_06814_),
    .B(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__a21o_1 _13974_ (.A1(_06804_),
    .A2(_06811_),
    .B1(_06809_),
    .X(_06817_));
 sky130_fd_sc_hd__xor2_1 _13975_ (.A(_06816_),
    .B(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__or2_1 _13976_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(_06819_));
 sky130_fd_sc_hd__o211a_1 _13977_ (.A1(_06555_),
    .A2(_06818_),
    .B1(_06819_),
    .C1(_06747_),
    .X(_00921_));
 sky130_fd_sc_hd__or2_1 _13978_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_06807_),
    .X(_06820_));
 sky130_fd_sc_hd__nand2_1 _13979_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_06807_),
    .Y(_06821_));
 sky130_fd_sc_hd__nand2_1 _13980_ (.A(_06820_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__a21o_1 _13981_ (.A1(_06815_),
    .A2(_06817_),
    .B1(_06814_),
    .X(_06823_));
 sky130_fd_sc_hd__xnor2_1 _13982_ (.A(_06822_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__mux2_1 _13983_ (.A0(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A1(_06824_),
    .S(_06553_),
    .X(_06825_));
 sky130_fd_sc_hd__and2_1 _13984_ (.A(_01253_),
    .B(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__clkbuf_1 _13985_ (.A(_06826_),
    .X(_00922_));
 sky130_fd_sc_hd__or2_1 _13986_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_06807_),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_1 _13987_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_06807_),
    .Y(_06828_));
 sky130_fd_sc_hd__nand2_1 _13988_ (.A(_06827_),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__a21bo_1 _13989_ (.A1(_06820_),
    .A2(_06823_),
    .B1_N(_06821_),
    .X(_06830_));
 sky130_fd_sc_hd__xnor2_1 _13990_ (.A(_06829_),
    .B(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__or2_1 _13991_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(_06832_));
 sky130_fd_sc_hd__o211a_1 _13992_ (.A1(_06555_),
    .A2(_06831_),
    .B1(_06832_),
    .C1(_06747_),
    .X(_00923_));
 sky130_fd_sc_hd__o21ai_1 _13993_ (.A1(_06809_),
    .A2(_06814_),
    .B1(_06815_),
    .Y(_06833_));
 sky130_fd_sc_hd__o311a_1 _13994_ (.A1(_06822_),
    .A2(_06833_),
    .A3(_06829_),
    .B1(_06828_),
    .C1(_06821_),
    .X(_06834_));
 sky130_fd_sc_hd__nand2_1 _13995_ (.A(_06811_),
    .B(_06816_),
    .Y(_06835_));
 sky130_fd_sc_hd__or4b_1 _13996_ (.A(_06822_),
    .B(_06835_),
    .C(_06829_),
    .D_N(_06804_),
    .X(_06836_));
 sky130_fd_sc_hd__buf_2 _13997_ (.A(_06807_),
    .X(_06837_));
 sky130_fd_sc_hd__xor2_1 _13998_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__a21boi_2 _13999_ (.A1(_06834_),
    .A2(_06836_),
    .B1_N(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__and3b_1 _14000_ (.A_N(_06838_),
    .B(_06834_),
    .C(_06836_),
    .X(_06840_));
 sky130_fd_sc_hd__o21ai_1 _14001_ (.A1(_06839_),
    .A2(_06840_),
    .B1(_06584_),
    .Y(_06841_));
 sky130_fd_sc_hd__o211a_1 _14002_ (.A1(_06561_),
    .A2(net462),
    .B1(_06678_),
    .C1(_06841_),
    .X(_00924_));
 sky130_fd_sc_hd__or2_1 _14003_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_06807_),
    .X(_06842_));
 sky130_fd_sc_hd__nand2_1 _14004_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_06837_),
    .Y(_06843_));
 sky130_fd_sc_hd__and2_1 _14005_ (.A(_06842_),
    .B(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__buf_2 _14006_ (.A(_06837_),
    .X(_06845_));
 sky130_fd_sc_hd__a21oi_1 _14007_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_06845_),
    .B1(_06839_),
    .Y(_06846_));
 sky130_fd_sc_hd__xnor2_1 _14008_ (.A(_06844_),
    .B(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__or2_1 _14009_ (.A(_06732_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_06848_));
 sky130_fd_sc_hd__o211a_1 _14010_ (.A1(_06555_),
    .A2(_06847_),
    .B1(_06848_),
    .C1(_06747_),
    .X(_00925_));
 sky130_fd_sc_hd__or2_1 _14011_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_06837_),
    .X(_06849_));
 sky130_fd_sc_hd__nand2_1 _14012_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_06837_),
    .Y(_06850_));
 sky130_fd_sc_hd__and2_1 _14013_ (.A(_06849_),
    .B(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__o21a_1 _14014_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_06845_),
    .X(_06852_));
 sky130_fd_sc_hd__a21oi_1 _14015_ (.A1(_06839_),
    .A2(_06842_),
    .B1(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__xnor2_1 _14016_ (.A(_06851_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__mux2_1 _14017_ (.A0(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A1(_06854_),
    .S(_06553_),
    .X(_06855_));
 sky130_fd_sc_hd__and2_1 _14018_ (.A(_01253_),
    .B(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__clkbuf_1 _14019_ (.A(_06856_),
    .X(_00926_));
 sky130_fd_sc_hd__or2b_1 _14020_ (.A(_06853_),
    .B_N(_06851_),
    .X(_06857_));
 sky130_fd_sc_hd__xor2_1 _14021_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_06837_),
    .X(_06858_));
 sky130_fd_sc_hd__a21oi_1 _14022_ (.A1(_06850_),
    .A2(_06857_),
    .B1(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__a31o_1 _14023_ (.A1(_06850_),
    .A2(_06857_),
    .A3(_06858_),
    .B1(_06569_),
    .X(_06860_));
 sky130_fd_sc_hd__o221a_1 _14024_ (.A1(_06563_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B1(_06859_),
    .B2(_06860_),
    .C1(_06631_),
    .X(_00927_));
 sky130_fd_sc_hd__or2_1 _14025_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_06837_),
    .X(_06861_));
 sky130_fd_sc_hd__nand2_1 _14026_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_06837_),
    .Y(_06862_));
 sky130_fd_sc_hd__and2_1 _14027_ (.A(_06861_),
    .B(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__and3_1 _14028_ (.A(_06844_),
    .B(_06851_),
    .C(_06858_),
    .X(_06864_));
 sky130_fd_sc_hd__o41a_1 _14029_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A4(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_06845_),
    .X(_06865_));
 sky130_fd_sc_hd__a21oi_2 _14030_ (.A1(_06839_),
    .A2(_06864_),
    .B1(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__xnor2_1 _14031_ (.A(_06863_),
    .B(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__or2_1 _14032_ (.A(_06562_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_06868_));
 sky130_fd_sc_hd__o211a_1 _14033_ (.A1(_06555_),
    .A2(_06867_),
    .B1(_06868_),
    .C1(_06747_),
    .X(_00928_));
 sky130_fd_sc_hd__or2b_1 _14034_ (.A(_06866_),
    .B_N(_06863_),
    .X(_06869_));
 sky130_fd_sc_hd__or2_1 _14035_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_06837_),
    .X(_06870_));
 sky130_fd_sc_hd__nand2_1 _14036_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_06837_),
    .Y(_06871_));
 sky130_fd_sc_hd__and2_1 _14037_ (.A(_06870_),
    .B(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__a21oi_1 _14038_ (.A1(_06862_),
    .A2(_06869_),
    .B1(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__a31o_1 _14039_ (.A1(_06862_),
    .A2(_06869_),
    .A3(_06872_),
    .B1(_06569_),
    .X(_06874_));
 sky130_fd_sc_hd__o221a_1 _14040_ (.A1(_06563_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_06873_),
    .B2(_06874_),
    .C1(_06631_),
    .X(_00929_));
 sky130_fd_sc_hd__inv_2 _14041_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .Y(_06875_));
 sky130_fd_sc_hd__or2_1 _14042_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06845_),
    .X(_06876_));
 sky130_fd_sc_hd__nand2_1 _14043_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_06845_),
    .Y(_06877_));
 sky130_fd_sc_hd__nand2_1 _14044_ (.A(_06876_),
    .B(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__nand2_1 _14045_ (.A(_06863_),
    .B(_06872_),
    .Y(_06879_));
 sky130_fd_sc_hd__o211a_1 _14046_ (.A1(_06866_),
    .A2(_06879_),
    .B1(_06871_),
    .C1(_06862_),
    .X(_06880_));
 sky130_fd_sc_hd__xnor2_1 _14047_ (.A(_06878_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__mux2_1 _14048_ (.A0(_06875_),
    .A1(_06881_),
    .S(_06562_),
    .X(_06882_));
 sky130_fd_sc_hd__and2b_1 _14049_ (.A_N(_06882_),
    .B(_01512_),
    .X(_06883_));
 sky130_fd_sc_hd__clkbuf_1 _14050_ (.A(_06883_),
    .X(_00930_));
 sky130_fd_sc_hd__or2_1 _14051_ (.A(_06878_),
    .B(_06880_),
    .X(_06884_));
 sky130_fd_sc_hd__xor2_1 _14052_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_06845_),
    .X(_06885_));
 sky130_fd_sc_hd__a21oi_1 _14053_ (.A1(_06877_),
    .A2(_06884_),
    .B1(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__a31o_1 _14054_ (.A1(_06877_),
    .A2(_06884_),
    .A3(_06885_),
    .B1(_06569_),
    .X(_06887_));
 sky130_fd_sc_hd__o221a_1 _14055_ (.A1(_06563_),
    .A2(net605),
    .B1(_06886_),
    .B2(_06887_),
    .C1(_06631_),
    .X(_00931_));
 sky130_fd_sc_hd__and2_1 _14056_ (.A(_06569_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .X(_06888_));
 sky130_fd_sc_hd__nor2_1 _14057_ (.A(_06878_),
    .B(_06879_),
    .Y(_06889_));
 sky130_fd_sc_hd__and4_1 _14058_ (.A(_06839_),
    .B(_06864_),
    .C(_06885_),
    .D(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__o41a_1 _14059_ (.A1(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .A3(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A4(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_06845_),
    .X(_06891_));
 sky130_fd_sc_hd__or2_1 _14060_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06845_),
    .X(_06892_));
 sky130_fd_sc_hd__nand2_1 _14061_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_06845_),
    .Y(_06893_));
 sky130_fd_sc_hd__and2_1 _14062_ (.A(_06892_),
    .B(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__o31ai_2 _14063_ (.A1(_06865_),
    .A2(_06890_),
    .A3(_06891_),
    .B1(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__or4_1 _14064_ (.A(_06865_),
    .B(_06894_),
    .C(_06890_),
    .D(_06891_),
    .X(_06896_));
 sky130_fd_sc_hd__and3_1 _14065_ (.A(_06557_),
    .B(_06895_),
    .C(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__o21a_1 _14066_ (.A1(_06888_),
    .A2(_06897_),
    .B1(_04961_),
    .X(_00932_));
 sky130_fd_sc_hd__xor2_1 _14067_ (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_06845_),
    .X(_06898_));
 sky130_fd_sc_hd__a21oi_1 _14068_ (.A1(_06893_),
    .A2(_06895_),
    .B1(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__a31o_1 _14069_ (.A1(_06893_),
    .A2(_06895_),
    .A3(_06898_),
    .B1(_06569_),
    .X(_06900_));
 sky130_fd_sc_hd__o221a_1 _14070_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .A2(_06565_),
    .B1(_06899_),
    .B2(_06900_),
    .C1(_06631_),
    .X(_00933_));
 sky130_fd_sc_hd__and2_1 _14071_ (.A(_06557_),
    .B(_01979_),
    .X(_06901_));
 sky130_fd_sc_hd__clkbuf_1 _14072_ (.A(_06901_),
    .X(_00934_));
 sky130_fd_sc_hd__inv_2 _14073_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.valid_out ),
    .Y(_06902_));
 sky130_fd_sc_hd__clkbuf_4 _14074_ (.A(_06902_),
    .X(_06903_));
 sky130_fd_sc_hd__clkbuf_4 _14075_ (.A(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__clkbuf_4 _14076_ (.A(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__or2_1 _14077_ (.A(_01862_),
    .B(_01010_),
    .X(_06906_));
 sky130_fd_sc_hd__o211a_1 _14078_ (.A1(_06905_),
    .A2(net256),
    .B1(_06678_),
    .C1(_06906_),
    .X(_00935_));
 sky130_fd_sc_hd__clkbuf_4 _14079_ (.A(_01861_),
    .X(_06907_));
 sky130_fd_sc_hd__or2_1 _14080_ (.A(_06907_),
    .B(_01022_),
    .X(_06908_));
 sky130_fd_sc_hd__o211a_1 _14081_ (.A1(_06905_),
    .A2(net263),
    .B1(_06678_),
    .C1(_06908_),
    .X(_00936_));
 sky130_fd_sc_hd__buf_2 _14082_ (.A(_01861_),
    .X(_06909_));
 sky130_fd_sc_hd__buf_4 _14083_ (.A(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__clkbuf_4 _14084_ (.A(_06909_),
    .X(_06911_));
 sky130_fd_sc_hd__nand2_1 _14085_ (.A(_06911_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .Y(_06912_));
 sky130_fd_sc_hd__o211a_1 _14086_ (.A1(_06910_),
    .A2(net245),
    .B1(_06678_),
    .C1(_06912_),
    .X(_00937_));
 sky130_fd_sc_hd__nand2_1 _14087_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .Y(_06913_));
 sky130_fd_sc_hd__or2_1 _14088_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_06914_));
 sky130_fd_sc_hd__a21oi_1 _14089_ (.A1(_06913_),
    .A2(_06914_),
    .B1(_06647_),
    .Y(_06915_));
 sky130_fd_sc_hd__a31o_1 _14090_ (.A1(_06647_),
    .A2(_06913_),
    .A3(_06914_),
    .B1(_06904_),
    .X(_06916_));
 sky130_fd_sc_hd__o221a_1 _14091_ (.A1(_06910_),
    .A2(net318),
    .B1(_06915_),
    .B2(_06916_),
    .C1(_06631_),
    .X(_00938_));
 sky130_fd_sc_hd__and3_1 _14092_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .C(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(_06917_));
 sky130_fd_sc_hd__a21oi_1 _14093_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .B1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .Y(_06918_));
 sky130_fd_sc_hd__or2_1 _14094_ (.A(_06917_),
    .B(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__nor2_1 _14095_ (.A(_06915_),
    .B(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__a21o_1 _14096_ (.A1(_06915_),
    .A2(_06919_),
    .B1(_06904_),
    .X(_06921_));
 sky130_fd_sc_hd__clkbuf_4 _14097_ (.A(_01474_),
    .X(_06922_));
 sky130_fd_sc_hd__o221a_1 _14098_ (.A1(_06910_),
    .A2(net323),
    .B1(_06920_),
    .B2(_06921_),
    .C1(_06922_),
    .X(_00939_));
 sky130_fd_sc_hd__nand2_1 _14099_ (.A(_06647_),
    .B(_06917_),
    .Y(_06923_));
 sky130_fd_sc_hd__or3_1 _14100_ (.A(_06646_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .C(_06914_),
    .X(_06924_));
 sky130_fd_sc_hd__a21oi_1 _14101_ (.A1(_06923_),
    .A2(_06924_),
    .B1(net358),
    .Y(_06925_));
 sky130_fd_sc_hd__clkbuf_4 _14102_ (.A(_06902_),
    .X(_06926_));
 sky130_fd_sc_hd__a31o_1 _14103_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A2(_06923_),
    .A3(_06924_),
    .B1(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__o221a_1 _14104_ (.A1(_06910_),
    .A2(net303),
    .B1(_06925_),
    .B2(_06927_),
    .C1(_06922_),
    .X(_00940_));
 sky130_fd_sc_hd__clkbuf_4 _14105_ (.A(_06909_),
    .X(_06928_));
 sky130_fd_sc_hd__or3_1 _14106_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .C(_06914_),
    .X(_06929_));
 sky130_fd_sc_hd__nand2_1 _14107_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .B(_06917_),
    .Y(_06930_));
 sky130_fd_sc_hd__mux2_1 _14108_ (.A0(_06929_),
    .A1(_06930_),
    .S(_06646_),
    .X(_06931_));
 sky130_fd_sc_hd__and2_1 _14109_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .B(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__o21ai_1 _14110_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_06931_),
    .B1(_01862_),
    .Y(_06933_));
 sky130_fd_sc_hd__o221a_1 _14111_ (.A1(_06928_),
    .A2(net316),
    .B1(_06932_),
    .B2(_06933_),
    .C1(_06922_),
    .X(_00941_));
 sky130_fd_sc_hd__inv_2 _14112_ (.A(_06646_),
    .Y(_06934_));
 sky130_fd_sc_hd__o21ai_1 _14113_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(_06929_),
    .B1(_06934_),
    .Y(_06935_));
 sky130_fd_sc_hd__a31o_1 _14114_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .A3(_06917_),
    .B1(_06934_),
    .X(_06936_));
 sky130_fd_sc_hd__inv_2 _14115_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .Y(_06937_));
 sky130_fd_sc_hd__a21oi_1 _14116_ (.A1(_06935_),
    .A2(_06936_),
    .B1(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__a31o_1 _14117_ (.A1(_06937_),
    .A2(_06935_),
    .A3(_06936_),
    .B1(_06926_),
    .X(_06939_));
 sky130_fd_sc_hd__o221a_1 _14118_ (.A1(_06928_),
    .A2(net339),
    .B1(_06938_),
    .B2(_06939_),
    .C1(_06922_),
    .X(_00942_));
 sky130_fd_sc_hd__and4_1 _14119_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .D(_06917_),
    .X(_06940_));
 sky130_fd_sc_hd__or3_1 _14120_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .C(_06929_),
    .X(_06941_));
 sky130_fd_sc_hd__inv_2 _14121_ (.A(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__mux2_1 _14122_ (.A0(_06940_),
    .A1(_06942_),
    .S(_06934_),
    .X(_06943_));
 sky130_fd_sc_hd__xnor2_1 _14123_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_1 _14124_ (.A(_06911_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__o211a_1 _14125_ (.A1(_06910_),
    .A2(net215),
    .B1(_06678_),
    .C1(_06945_),
    .X(_00943_));
 sky130_fd_sc_hd__or2_1 _14126_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .B(_06941_),
    .X(_06946_));
 sky130_fd_sc_hd__nor2_1 _14127_ (.A(_06646_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__a31o_1 _14128_ (.A1(_06647_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .A3(_06940_),
    .B1(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__xor2_1 _14129_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__or2_1 _14130_ (.A(_06907_),
    .B(net348),
    .X(_06950_));
 sky130_fd_sc_hd__o211a_1 _14131_ (.A1(_06905_),
    .A2(_06949_),
    .B1(_06950_),
    .C1(_06747_),
    .X(_00944_));
 sky130_fd_sc_hd__and3_1 _14132_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .C(_06940_),
    .X(_06951_));
 sky130_fd_sc_hd__nand2_1 _14133_ (.A(_06646_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__o31a_1 _14134_ (.A1(_06647_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A3(_06946_),
    .B1(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__and2_1 _14135_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .B(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__o21ai_1 _14136_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A2(_06953_),
    .B1(_01862_),
    .Y(_06955_));
 sky130_fd_sc_hd__o221a_1 _14137_ (.A1(_06928_),
    .A2(net334),
    .B1(_06954_),
    .B2(_06955_),
    .C1(_06922_),
    .X(_00945_));
 sky130_fd_sc_hd__nand3_1 _14138_ (.A(_06647_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(_06951_),
    .Y(_06956_));
 sky130_fd_sc_hd__o41a_1 _14139_ (.A1(_06646_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .A3(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .A4(_06946_),
    .B1(_06956_),
    .X(_06957_));
 sky130_fd_sc_hd__nor2_1 _14140_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__a21o_1 _14141_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .A2(_06957_),
    .B1(_06904_),
    .X(_06959_));
 sky130_fd_sc_hd__o221a_1 _14142_ (.A1(_06928_),
    .A2(net346),
    .B1(_06958_),
    .B2(_06959_),
    .C1(_06922_),
    .X(_00946_));
 sky130_fd_sc_hd__or4_1 _14143_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .D(_06946_),
    .X(_06960_));
 sky130_fd_sc_hd__and3_1 _14144_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .C(_06951_),
    .X(_06961_));
 sky130_fd_sc_hd__nand2_1 _14145_ (.A(_06646_),
    .B(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__o21a_1 _14146_ (.A1(_06647_),
    .A2(_06960_),
    .B1(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__and2_1 _14147_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__o21ai_1 _14148_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .A2(_06963_),
    .B1(_01862_),
    .Y(_06965_));
 sky130_fd_sc_hd__o221a_1 _14149_ (.A1(_06928_),
    .A2(net322),
    .B1(_06964_),
    .B2(_06965_),
    .C1(_06922_),
    .X(_00947_));
 sky130_fd_sc_hd__inv_2 _14150_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .Y(_06966_));
 sky130_fd_sc_hd__and2_1 _14151_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_06961_),
    .X(_06967_));
 sky130_fd_sc_hd__nor2_1 _14152_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .B(_06960_),
    .Y(_06968_));
 sky130_fd_sc_hd__mux2_1 _14153_ (.A0(_06967_),
    .A1(_06968_),
    .S(_06934_),
    .X(_06969_));
 sky130_fd_sc_hd__a21oi_1 _14154_ (.A1(_06966_),
    .A2(_06969_),
    .B1(_06904_),
    .Y(_06970_));
 sky130_fd_sc_hd__o21ai_1 _14155_ (.A1(_06966_),
    .A2(_06969_),
    .B1(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__o211a_1 _14156_ (.A1(_06910_),
    .A2(net236),
    .B1(_06678_),
    .C1(_06971_),
    .X(_00948_));
 sky130_fd_sc_hd__nand2_1 _14157_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .B(_06967_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand2_1 _14158_ (.A(_06966_),
    .B(_06968_),
    .Y(_06973_));
 sky130_fd_sc_hd__mux2_1 _14159_ (.A0(_06972_),
    .A1(_06973_),
    .S(_06934_),
    .X(_06974_));
 sky130_fd_sc_hd__nor2_1 _14160_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__a21o_1 _14161_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .A2(_06974_),
    .B1(_06904_),
    .X(_06976_));
 sky130_fd_sc_hd__o221a_1 _14162_ (.A1(_06928_),
    .A2(net320),
    .B1(_06975_),
    .B2(_06976_),
    .C1(_06922_),
    .X(_00949_));
 sky130_fd_sc_hd__or2_1 _14163_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(_06973_),
    .X(_06977_));
 sky130_fd_sc_hd__and3_1 _14164_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .C(_06967_),
    .X(_06978_));
 sky130_fd_sc_hd__nand2_1 _14165_ (.A(_06646_),
    .B(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__o21a_1 _14166_ (.A1(_06647_),
    .A2(_06977_),
    .B1(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__and2_1 _14167_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__o21ai_1 _14168_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A2(_06980_),
    .B1(_01862_),
    .Y(_06982_));
 sky130_fd_sc_hd__o221a_1 _14169_ (.A1(_06928_),
    .A2(net317),
    .B1(_06981_),
    .B2(_06982_),
    .C1(_06922_),
    .X(_00950_));
 sky130_fd_sc_hd__nand2_1 _14170_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_06978_),
    .Y(_06983_));
 sky130_fd_sc_hd__or2_1 _14171_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .B(_06977_),
    .X(_06984_));
 sky130_fd_sc_hd__mux2_1 _14172_ (.A0(_06983_),
    .A1(_06984_),
    .S(_06934_),
    .X(_06985_));
 sky130_fd_sc_hd__and2_1 _14173_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .B(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__o21ai_1 _14174_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A2(_06985_),
    .B1(_01862_),
    .Y(_06987_));
 sky130_fd_sc_hd__o221a_1 _14175_ (.A1(_06928_),
    .A2(net278),
    .B1(_06986_),
    .B2(_06987_),
    .C1(_06922_),
    .X(_00951_));
 sky130_fd_sc_hd__xor2_1 _14176_ (.A(_06647_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(_06988_));
 sky130_fd_sc_hd__o21a_1 _14177_ (.A1(_06985_),
    .A2(_06988_),
    .B1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(_06989_));
 sky130_fd_sc_hd__o31ai_1 _14178_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(_06985_),
    .A3(_06988_),
    .B1(_01862_),
    .Y(_06990_));
 sky130_fd_sc_hd__o221a_1 _14179_ (.A1(_06928_),
    .A2(net293),
    .B1(_06989_),
    .B2(_06990_),
    .C1(_01456_),
    .X(_00952_));
 sky130_fd_sc_hd__o31a_1 _14180_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(_06984_),
    .B1(_06934_),
    .X(_06991_));
 sky130_fd_sc_hd__a41o_1 _14181_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .A3(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .A4(_06978_),
    .B1(_06934_),
    .X(_06992_));
 sky130_fd_sc_hd__or2b_1 _14182_ (.A(_06991_),
    .B_N(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__xnor2_1 _14183_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .B(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__or2_1 _14184_ (.A(_06907_),
    .B(net432),
    .X(_06995_));
 sky130_fd_sc_hd__clkbuf_4 _14185_ (.A(_04455_),
    .X(_06996_));
 sky130_fd_sc_hd__o211a_1 _14186_ (.A1(_06905_),
    .A2(_06994_),
    .B1(_06995_),
    .C1(_06996_),
    .X(_00953_));
 sky130_fd_sc_hd__a21oi_1 _14187_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .A2(_06992_),
    .B1(_06991_),
    .Y(_06997_));
 sky130_fd_sc_hd__or2_1 _14188_ (.A(_06907_),
    .B(net412),
    .X(_06998_));
 sky130_fd_sc_hd__o211a_1 _14189_ (.A1(_06905_),
    .A2(_06997_),
    .B1(_06998_),
    .C1(_06996_),
    .X(_00954_));
 sky130_fd_sc_hd__nor2_1 _14190_ (.A(_06875_),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .Y(_06999_));
 sky130_fd_sc_hd__a21o_1 _14191_ (.A1(_06875_),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_06904_),
    .X(_07000_));
 sky130_fd_sc_hd__o221a_1 _14192_ (.A1(_06928_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .B1(_06999_),
    .B2(_07000_),
    .C1(_01456_),
    .X(_00955_));
 sky130_fd_sc_hd__and2b_1 _14193_ (.A_N(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_07001_));
 sky130_fd_sc_hd__xnor2_2 _14194_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__xnor2_2 _14195_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__xor2_1 _14196_ (.A(_06999_),
    .B(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__or2_1 _14197_ (.A(_06907_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(_07005_));
 sky130_fd_sc_hd__o211a_1 _14198_ (.A1(_06905_),
    .A2(_07004_),
    .B1(_07005_),
    .C1(_06996_),
    .X(_00956_));
 sky130_fd_sc_hd__o21ba_1 _14199_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B1_N(_06646_),
    .X(_07006_));
 sky130_fd_sc_hd__xnor2_1 _14200_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__nor2_1 _14201_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__and2_1 _14202_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B(_07007_),
    .X(_07009_));
 sky130_fd_sc_hd__nor2_1 _14203_ (.A(_07008_),
    .B(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__nand2_1 _14204_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .B(_07002_),
    .Y(_07011_));
 sky130_fd_sc_hd__o21ai_2 _14205_ (.A1(_06999_),
    .A2(_07003_),
    .B1(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__nand2_1 _14206_ (.A(_07010_),
    .B(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__o21a_1 _14207_ (.A1(_07010_),
    .A2(_07012_),
    .B1(_01861_),
    .X(_07014_));
 sky130_fd_sc_hd__a22o_1 _14208_ (.A1(_06903_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ),
    .B1(_07013_),
    .B2(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__and2_1 _14209_ (.A(_01253_),
    .B(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__clkbuf_1 _14210_ (.A(_07016_),
    .X(_00957_));
 sky130_fd_sc_hd__and2_1 _14211_ (.A(_06904_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .X(_07017_));
 sky130_fd_sc_hd__or2_1 _14212_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(_07018_));
 sky130_fd_sc_hd__or3b_1 _14213_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_07018_),
    .C_N(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_07019_));
 sky130_fd_sc_hd__o21ai_1 _14214_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_07018_),
    .B1(_06934_),
    .Y(_07020_));
 sky130_fd_sc_hd__mux2_1 _14215_ (.A0(_07020_),
    .A1(_06934_),
    .S(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(_07021_));
 sky130_fd_sc_hd__and3_1 _14216_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .B(_07019_),
    .C(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__clkbuf_4 _14217_ (.A(_07021_),
    .X(_07023_));
 sky130_fd_sc_hd__a21oi_1 _14218_ (.A1(_07019_),
    .A2(_07023_),
    .B1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[3] ),
    .Y(_07024_));
 sky130_fd_sc_hd__or2_1 _14219_ (.A(_07022_),
    .B(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__a21oi_1 _14220_ (.A1(_07010_),
    .A2(_07012_),
    .B1(_07009_),
    .Y(_07026_));
 sky130_fd_sc_hd__o21ai_1 _14221_ (.A1(_07025_),
    .A2(_07026_),
    .B1(_01862_),
    .Y(_07027_));
 sky130_fd_sc_hd__a21oi_1 _14222_ (.A1(_07025_),
    .A2(_07026_),
    .B1(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__o21a_1 _14223_ (.A1(_07017_),
    .A2(_07028_),
    .B1(_04961_),
    .X(_00958_));
 sky130_fd_sc_hd__o21ba_1 _14224_ (.A1(_07024_),
    .A2(_07026_),
    .B1_N(_07022_),
    .X(_07029_));
 sky130_fd_sc_hd__nand2_1 _14225_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_07023_),
    .Y(_07030_));
 sky130_fd_sc_hd__or2_1 _14226_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B(_07021_),
    .X(_07031_));
 sky130_fd_sc_hd__nand2_1 _14227_ (.A(_07030_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__xor2_1 _14228_ (.A(_07029_),
    .B(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__or2_1 _14229_ (.A(_06907_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(_07034_));
 sky130_fd_sc_hd__o211a_1 _14230_ (.A1(_06905_),
    .A2(_07033_),
    .B1(_07034_),
    .C1(_06996_),
    .X(_00959_));
 sky130_fd_sc_hd__xnor2_1 _14231_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .B(_07023_),
    .Y(_07035_));
 sky130_fd_sc_hd__o21ai_1 _14232_ (.A1(_07029_),
    .A2(_07032_),
    .B1(_07030_),
    .Y(_07036_));
 sky130_fd_sc_hd__xnor2_1 _14233_ (.A(_07035_),
    .B(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__or2_1 _14234_ (.A(_06907_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(_07038_));
 sky130_fd_sc_hd__o211a_1 _14235_ (.A1(_06905_),
    .A2(_07037_),
    .B1(_07038_),
    .C1(_06996_),
    .X(_00960_));
 sky130_fd_sc_hd__nor2_1 _14236_ (.A(_07032_),
    .B(_07035_),
    .Y(_07039_));
 sky130_fd_sc_hd__and2b_1 _14237_ (.A_N(_07029_),
    .B(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__buf_4 _14238_ (.A(_07023_),
    .X(_07041_));
 sky130_fd_sc_hd__clkbuf_4 _14239_ (.A(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__o21a_1 _14240_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B1(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__nand2_1 _14241_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_07023_),
    .Y(_07044_));
 sky130_fd_sc_hd__or2_1 _14242_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B(_07023_),
    .X(_07045_));
 sky130_fd_sc_hd__and2_1 _14243_ (.A(_07044_),
    .B(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__o21ai_1 _14244_ (.A1(_07040_),
    .A2(_07043_),
    .B1(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__o31a_1 _14245_ (.A1(_07046_),
    .A2(_07040_),
    .A3(_07043_),
    .B1(_01861_),
    .X(_07048_));
 sky130_fd_sc_hd__a22oi_1 _14246_ (.A1(_06903_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .B1(_07047_),
    .B2(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__and2b_1 _14247_ (.A_N(_07049_),
    .B(_01512_),
    .X(_07050_));
 sky130_fd_sc_hd__clkbuf_1 _14248_ (.A(_07050_),
    .X(_00961_));
 sky130_fd_sc_hd__xor2_1 _14249_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B(_07023_),
    .X(_07051_));
 sky130_fd_sc_hd__a21oi_1 _14250_ (.A1(_07044_),
    .A2(_07047_),
    .B1(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__a31o_1 _14251_ (.A1(_07044_),
    .A2(_07047_),
    .A3(_07051_),
    .B1(_06926_),
    .X(_07053_));
 sky130_fd_sc_hd__o221a_1 _14252_ (.A1(_06911_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .B1(_07052_),
    .B2(_07053_),
    .C1(_01456_),
    .X(_00962_));
 sky130_fd_sc_hd__and4b_1 _14253_ (.A_N(_07029_),
    .B(_07046_),
    .C(_07039_),
    .D(_07051_),
    .X(_07054_));
 sky130_fd_sc_hd__o41a_1 _14254_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .A3(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .A4(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .B1(_07041_),
    .X(_07055_));
 sky130_fd_sc_hd__xor2_1 _14255_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B(_07041_),
    .X(_07056_));
 sky130_fd_sc_hd__o21ai_2 _14256_ (.A1(_07054_),
    .A2(_07055_),
    .B1(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__or3_1 _14257_ (.A(_07056_),
    .B(_07054_),
    .C(_07055_),
    .X(_07058_));
 sky130_fd_sc_hd__clkbuf_4 _14258_ (.A(_06903_),
    .X(_07059_));
 sky130_fd_sc_hd__a21o_1 _14259_ (.A1(_07057_),
    .A2(_07058_),
    .B1(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__o211a_1 _14260_ (.A1(_06910_),
    .A2(net587),
    .B1(_06678_),
    .C1(_07060_),
    .X(_00963_));
 sky130_fd_sc_hd__xnor2_1 _14261_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .B(_07023_),
    .Y(_07061_));
 sky130_fd_sc_hd__a21bo_1 _14262_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .A2(_07042_),
    .B1_N(_07057_),
    .X(_07062_));
 sky130_fd_sc_hd__xnor2_1 _14263_ (.A(_07061_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__or2_1 _14264_ (.A(_06907_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(_07064_));
 sky130_fd_sc_hd__o211a_1 _14265_ (.A1(_06905_),
    .A2(_07063_),
    .B1(_07064_),
    .C1(_06996_),
    .X(_00964_));
 sky130_fd_sc_hd__o21bai_1 _14266_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(_07042_),
    .B1_N(_07057_),
    .Y(_07065_));
 sky130_fd_sc_hd__o21ai_1 _14267_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_07042_),
    .Y(_07066_));
 sky130_fd_sc_hd__xnor2_1 _14268_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B(_07041_),
    .Y(_07067_));
 sky130_fd_sc_hd__a21oi_1 _14269_ (.A1(_07065_),
    .A2(_07066_),
    .B1(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__a31o_1 _14270_ (.A1(_07067_),
    .A2(_07065_),
    .A3(_07066_),
    .B1(_06902_),
    .X(_07069_));
 sky130_fd_sc_hd__o2bb2a_1 _14271_ (.A1_N(_06903_),
    .A2_N(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .B1(_07068_),
    .B2(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__and2b_1 _14272_ (.A_N(_07070_),
    .B(_01512_),
    .X(_07071_));
 sky130_fd_sc_hd__clkbuf_1 _14273_ (.A(_07071_),
    .X(_00965_));
 sky130_fd_sc_hd__xnor2_1 _14274_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .B(_07041_),
    .Y(_07072_));
 sky130_fd_sc_hd__a21o_1 _14275_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A2(_07042_),
    .B1(_07068_),
    .X(_07073_));
 sky130_fd_sc_hd__xnor2_1 _14276_ (.A(_07072_),
    .B(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__or2_1 _14277_ (.A(_06907_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(_07075_));
 sky130_fd_sc_hd__o211a_1 _14278_ (.A1(_06905_),
    .A2(_07074_),
    .B1(_07075_),
    .C1(_06996_),
    .X(_00966_));
 sky130_fd_sc_hd__and2_1 _14279_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_07023_),
    .X(_07076_));
 sky130_fd_sc_hd__or2_1 _14280_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B(_07023_),
    .X(_07077_));
 sky130_fd_sc_hd__or2b_1 _14281_ (.A(_07076_),
    .B_N(_07077_),
    .X(_07078_));
 sky130_fd_sc_hd__or3_1 _14282_ (.A(_07061_),
    .B(_07067_),
    .C(_07072_),
    .X(_07079_));
 sky130_fd_sc_hd__o41ai_4 _14283_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .A3(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .A4(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .B1(_07041_),
    .Y(_07080_));
 sky130_fd_sc_hd__o21ai_2 _14284_ (.A1(_07057_),
    .A2(_07079_),
    .B1(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__xnor2_1 _14285_ (.A(_07078_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__or2_1 _14286_ (.A(_06907_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(_07083_));
 sky130_fd_sc_hd__o211a_1 _14287_ (.A1(_07059_),
    .A2(_07082_),
    .B1(_07083_),
    .C1(_06996_),
    .X(_00967_));
 sky130_fd_sc_hd__xnor2_1 _14288_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .B(_07041_),
    .Y(_07084_));
 sky130_fd_sc_hd__a21o_1 _14289_ (.A1(_07077_),
    .A2(_07081_),
    .B1(_07076_),
    .X(_07085_));
 sky130_fd_sc_hd__xnor2_1 _14290_ (.A(_07084_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__or2_1 _14291_ (.A(_06909_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(_07087_));
 sky130_fd_sc_hd__o211a_1 _14292_ (.A1(_07059_),
    .A2(_07086_),
    .B1(_07087_),
    .C1(_06996_),
    .X(_00968_));
 sky130_fd_sc_hd__xor2_1 _14293_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B(_07041_),
    .X(_07088_));
 sky130_fd_sc_hd__o21a_1 _14294_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .B1(_07041_),
    .X(_07089_));
 sky130_fd_sc_hd__nor2_1 _14295_ (.A(_07078_),
    .B(_07084_),
    .Y(_07090_));
 sky130_fd_sc_hd__and2_1 _14296_ (.A(_07081_),
    .B(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__o31ai_1 _14297_ (.A1(_07088_),
    .A2(_07089_),
    .A3(_07091_),
    .B1(_01861_),
    .Y(_07092_));
 sky130_fd_sc_hd__o21a_1 _14298_ (.A1(_07089_),
    .A2(_07091_),
    .B1(_07088_),
    .X(_07093_));
 sky130_fd_sc_hd__a2bb2o_1 _14299_ (.A1_N(_07092_),
    .A2_N(_07093_),
    .B1(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B2(_06903_),
    .X(_07094_));
 sky130_fd_sc_hd__and2_1 _14300_ (.A(_01253_),
    .B(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__clkbuf_1 _14301_ (.A(_07095_),
    .X(_00969_));
 sky130_fd_sc_hd__xnor2_1 _14302_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_07041_),
    .Y(_07096_));
 sky130_fd_sc_hd__a21o_1 _14303_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .A2(_07042_),
    .B1(_07093_),
    .X(_07097_));
 sky130_fd_sc_hd__xnor2_1 _14304_ (.A(_07096_),
    .B(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__or2_1 _14305_ (.A(_06909_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(_07099_));
 sky130_fd_sc_hd__o211a_1 _14306_ (.A1(_07059_),
    .A2(_07098_),
    .B1(_07099_),
    .C1(_06996_),
    .X(_00970_));
 sky130_fd_sc_hd__and2_1 _14307_ (.A(_06904_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .X(_07100_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(_07088_),
    .B(_07090_),
    .Y(_07101_));
 sky130_fd_sc_hd__or4_1 _14309_ (.A(_07057_),
    .B(_07079_),
    .C(_07096_),
    .D(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__o21a_1 _14310_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1(_07042_),
    .X(_07103_));
 sky130_fd_sc_hd__nor2_1 _14311_ (.A(_07089_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__xnor2_1 _14312_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_07042_),
    .Y(_07105_));
 sky130_fd_sc_hd__a31oi_1 _14313_ (.A1(_07080_),
    .A2(_07102_),
    .A3(_07104_),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__a41o_1 _14314_ (.A1(_07080_),
    .A2(_07105_),
    .A3(_07102_),
    .A4(_07104_),
    .B1(_06926_),
    .X(_07107_));
 sky130_fd_sc_hd__nor2_1 _14315_ (.A(_07106_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__o21a_1 _14316_ (.A1(_07100_),
    .A2(_07108_),
    .B1(_04961_),
    .X(_00971_));
 sky130_fd_sc_hd__a21o_1 _14317_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .A2(_07042_),
    .B1(_07106_),
    .X(_07109_));
 sky130_fd_sc_hd__xnor2_1 _14318_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .B(_07042_),
    .Y(_07110_));
 sky130_fd_sc_hd__xnor2_1 _14319_ (.A(_07109_),
    .B(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__or2_1 _14320_ (.A(_06909_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_07112_));
 sky130_fd_sc_hd__o211a_1 _14321_ (.A1(_07059_),
    .A2(_07111_),
    .B1(_07112_),
    .C1(_01475_),
    .X(_00972_));
 sky130_fd_sc_hd__and2_1 _14322_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .X(_07113_));
 sky130_fd_sc_hd__nor2_1 _14323_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .Y(_07114_));
 sky130_fd_sc_hd__o21ai_1 _14324_ (.A1(_07113_),
    .A2(_07114_),
    .B1(_06911_),
    .Y(_07115_));
 sky130_fd_sc_hd__o211a_1 _14325_ (.A1(_06910_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .B1(_01766_),
    .C1(_07115_),
    .X(_00973_));
 sky130_fd_sc_hd__and2b_1 _14326_ (.A_N(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .X(_07116_));
 sky130_fd_sc_hd__xnor2_1 _14327_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .B(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__xnor2_1 _14328_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .B(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__or2_1 _14329_ (.A(_07113_),
    .B(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__nand2_1 _14330_ (.A(_07113_),
    .B(_07118_),
    .Y(_07120_));
 sky130_fd_sc_hd__a21o_1 _14331_ (.A1(_07119_),
    .A2(_07120_),
    .B1(_06904_),
    .X(_07121_));
 sky130_fd_sc_hd__o211a_1 _14332_ (.A1(_06910_),
    .A2(net423),
    .B1(_01766_),
    .C1(_07121_),
    .X(_00974_));
 sky130_fd_sc_hd__nor2_1 _14333_ (.A(_01862_),
    .B(_01032_),
    .Y(_07122_));
 sky130_fd_sc_hd__or2b_1 _14334_ (.A(_07117_),
    .B_N(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(_07123_));
 sky130_fd_sc_hd__inv_2 _14335_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[2] ),
    .Y(_07124_));
 sky130_fd_sc_hd__o21ba_1 _14336_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .B1_N(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(_07125_));
 sky130_fd_sc_hd__xnor2_1 _14337_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__and2_1 _14338_ (.A(_07124_),
    .B(_07126_),
    .X(_07127_));
 sky130_fd_sc_hd__nor2_1 _14339_ (.A(_07124_),
    .B(_07126_),
    .Y(_07128_));
 sky130_fd_sc_hd__or2_1 _14340_ (.A(_07127_),
    .B(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__a21oi_1 _14341_ (.A1(_07123_),
    .A2(_07120_),
    .B1(_07129_),
    .Y(_07130_));
 sky130_fd_sc_hd__a31o_1 _14342_ (.A1(_07123_),
    .A2(_07120_),
    .A3(_07129_),
    .B1(_06926_),
    .X(_07131_));
 sky130_fd_sc_hd__nor2_1 _14343_ (.A(_07130_),
    .B(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__o21a_1 _14344_ (.A1(_07122_),
    .A2(_07132_),
    .B1(_01552_),
    .X(_00975_));
 sky130_fd_sc_hd__nor3_1 _14345_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ),
    .B(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .C(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ),
    .Y(_07133_));
 sky130_fd_sc_hd__nor2_1 _14346_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__mux2_1 _14347_ (.A0(_07134_),
    .A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .S(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(_07135_));
 sky130_fd_sc_hd__a21o_1 _14348_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .A2(_07133_),
    .B1(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__xor2_1 _14349_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__nor3_1 _14350_ (.A(_07128_),
    .B(_07130_),
    .C(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__o21a_1 _14351_ (.A1(_07128_),
    .A2(_07130_),
    .B1(_07137_),
    .X(_07139_));
 sky130_fd_sc_hd__nand2_1 _14352_ (.A(_06903_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .Y(_07140_));
 sky130_fd_sc_hd__o31ai_1 _14353_ (.A1(_06903_),
    .A2(_07138_),
    .A3(_07139_),
    .B1(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__and2_1 _14354_ (.A(_01253_),
    .B(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__clkbuf_1 _14355_ (.A(_07142_),
    .X(_00976_));
 sky130_fd_sc_hd__and2_1 _14356_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[3] ),
    .B(_07136_),
    .X(_07143_));
 sky130_fd_sc_hd__clkbuf_4 _14357_ (.A(_07135_),
    .X(_07144_));
 sky130_fd_sc_hd__or2_1 _14358_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B(_07144_),
    .Y(_07146_));
 sky130_fd_sc_hd__and2_1 _14360_ (.A(_07145_),
    .B(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__o21ai_1 _14361_ (.A1(_07143_),
    .A2(_07139_),
    .B1(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__or3_1 _14362_ (.A(_07143_),
    .B(_07139_),
    .C(_07147_),
    .X(_07149_));
 sky130_fd_sc_hd__and2_1 _14363_ (.A(_07148_),
    .B(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__or2_1 _14364_ (.A(_06909_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(_07151_));
 sky130_fd_sc_hd__o211a_1 _14365_ (.A1(_07059_),
    .A2(_07150_),
    .B1(_07151_),
    .C1(_01475_),
    .X(_00977_));
 sky130_fd_sc_hd__xor2_1 _14366_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .B(_07144_),
    .X(_07152_));
 sky130_fd_sc_hd__a21oi_1 _14367_ (.A1(_07146_),
    .A2(_07148_),
    .B1(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__a31o_1 _14368_ (.A1(_07146_),
    .A2(_07148_),
    .A3(_07152_),
    .B1(_06926_),
    .X(_07154_));
 sky130_fd_sc_hd__o221a_1 _14369_ (.A1(_06911_),
    .A2(net624),
    .B1(_07153_),
    .B2(_07154_),
    .C1(_01456_),
    .X(_00978_));
 sky130_fd_sc_hd__o211a_1 _14370_ (.A1(_07143_),
    .A2(_07139_),
    .B1(_07147_),
    .C1(_07152_),
    .X(_07155_));
 sky130_fd_sc_hd__clkbuf_4 _14371_ (.A(_07144_),
    .X(_07156_));
 sky130_fd_sc_hd__clkbuf_4 _14372_ (.A(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__o21a_1 _14373_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B1(_07157_),
    .X(_07158_));
 sky130_fd_sc_hd__or2_1 _14374_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_07144_),
    .X(_07159_));
 sky130_fd_sc_hd__nand2_1 _14375_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B(_07144_),
    .Y(_07160_));
 sky130_fd_sc_hd__and2_1 _14376_ (.A(_07159_),
    .B(_07160_),
    .X(_07161_));
 sky130_fd_sc_hd__o21ai_1 _14377_ (.A1(_07155_),
    .A2(_07158_),
    .B1(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__o31a_1 _14378_ (.A1(_07161_),
    .A2(_07155_),
    .A3(_07158_),
    .B1(_01861_),
    .X(_07163_));
 sky130_fd_sc_hd__a22o_1 _14379_ (.A1(_06903_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .B1(_07162_),
    .B2(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__and2_1 _14380_ (.A(_01253_),
    .B(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__clkbuf_1 _14381_ (.A(_07165_),
    .X(_00979_));
 sky130_fd_sc_hd__xor2_1 _14382_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B(_07144_),
    .X(_07166_));
 sky130_fd_sc_hd__a21oi_1 _14383_ (.A1(_07160_),
    .A2(_07162_),
    .B1(_07166_),
    .Y(_07167_));
 sky130_fd_sc_hd__a31o_1 _14384_ (.A1(_07160_),
    .A2(_07162_),
    .A3(_07166_),
    .B1(_06926_),
    .X(_07168_));
 sky130_fd_sc_hd__o221a_1 _14385_ (.A1(_06911_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .B1(_07167_),
    .B2(_07168_),
    .C1(_01456_),
    .X(_00980_));
 sky130_fd_sc_hd__and3_1 _14386_ (.A(_07161_),
    .B(_07155_),
    .C(_07166_),
    .X(_07169_));
 sky130_fd_sc_hd__o41a_1 _14387_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[6] ),
    .A3(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .A4(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .B1(_07156_),
    .X(_07170_));
 sky130_fd_sc_hd__xor2_1 _14388_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B(_07156_),
    .X(_07171_));
 sky130_fd_sc_hd__o21a_1 _14389_ (.A1(_07169_),
    .A2(_07170_),
    .B1(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__nor3_1 _14390_ (.A(_07171_),
    .B(_07169_),
    .C(_07170_),
    .Y(_07173_));
 sky130_fd_sc_hd__o21ai_1 _14391_ (.A1(_07172_),
    .A2(_07173_),
    .B1(_06911_),
    .Y(_07174_));
 sky130_fd_sc_hd__o211a_1 _14392_ (.A1(_06910_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_01766_),
    .C1(_07174_),
    .X(_00981_));
 sky130_fd_sc_hd__xor2_1 _14393_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .B(_07156_),
    .X(_07175_));
 sky130_fd_sc_hd__a21oi_1 _14394_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .A2(_07157_),
    .B1(_07172_),
    .Y(_07176_));
 sky130_fd_sc_hd__xnor2_1 _14395_ (.A(_07175_),
    .B(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__or2_1 _14396_ (.A(_06909_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(_07178_));
 sky130_fd_sc_hd__o211a_1 _14397_ (.A1(_07059_),
    .A2(_07177_),
    .B1(_07178_),
    .C1(_01475_),
    .X(_00982_));
 sky130_fd_sc_hd__o21a_1 _14398_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(_07157_),
    .B1(_07172_),
    .X(_07179_));
 sky130_fd_sc_hd__o21a_1 _14399_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_07157_),
    .X(_07180_));
 sky130_fd_sc_hd__or2_1 _14400_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_07144_),
    .X(_07181_));
 sky130_fd_sc_hd__nand2_1 _14401_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B(_07156_),
    .Y(_07182_));
 sky130_fd_sc_hd__and2_1 _14402_ (.A(_07181_),
    .B(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__o21ai_1 _14403_ (.A1(_07179_),
    .A2(_07180_),
    .B1(_07183_),
    .Y(_07184_));
 sky130_fd_sc_hd__o31a_1 _14404_ (.A1(_07183_),
    .A2(_07179_),
    .A3(_07180_),
    .B1(_01861_),
    .X(_07185_));
 sky130_fd_sc_hd__a22o_1 _14405_ (.A1(_06903_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .B1(_07184_),
    .B2(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__and2_1 _14406_ (.A(_01253_),
    .B(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__clkbuf_1 _14407_ (.A(_07187_),
    .X(_00983_));
 sky130_fd_sc_hd__xor2_1 _14408_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .B(_07156_),
    .X(_07188_));
 sky130_fd_sc_hd__a21oi_1 _14409_ (.A1(_07182_),
    .A2(_07184_),
    .B1(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__a31o_1 _14410_ (.A1(_07182_),
    .A2(_07184_),
    .A3(_07188_),
    .B1(_06926_),
    .X(_07190_));
 sky130_fd_sc_hd__o221a_1 _14411_ (.A1(_06911_),
    .A2(net549),
    .B1(_07189_),
    .B2(_07190_),
    .C1(_01456_),
    .X(_00984_));
 sky130_fd_sc_hd__or2_1 _14412_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_07144_),
    .X(_07191_));
 sky130_fd_sc_hd__nand2_1 _14413_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B(_07156_),
    .Y(_07192_));
 sky130_fd_sc_hd__and2_1 _14414_ (.A(_07191_),
    .B(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__and3_1 _14415_ (.A(_07175_),
    .B(_07183_),
    .C(_07188_),
    .X(_07194_));
 sky130_fd_sc_hd__o41a_1 _14416_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .A3(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .A4(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .B1(_07157_),
    .X(_07195_));
 sky130_fd_sc_hd__a21oi_1 _14417_ (.A1(_07172_),
    .A2(_07194_),
    .B1(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__xnor2_1 _14418_ (.A(_07193_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__or2_1 _14419_ (.A(_06909_),
    .B(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(_07198_));
 sky130_fd_sc_hd__o211a_1 _14420_ (.A1(_07059_),
    .A2(_07197_),
    .B1(_07198_),
    .C1(_01475_),
    .X(_00985_));
 sky130_fd_sc_hd__or2b_1 _14421_ (.A(_07196_),
    .B_N(_07193_),
    .X(_07199_));
 sky130_fd_sc_hd__xor2_1 _14422_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B(_07144_),
    .X(_07200_));
 sky130_fd_sc_hd__a21oi_1 _14423_ (.A1(_07192_),
    .A2(_07199_),
    .B1(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__a31o_1 _14424_ (.A1(_07192_),
    .A2(_07199_),
    .A3(_07200_),
    .B1(_06926_),
    .X(_07202_));
 sky130_fd_sc_hd__o221a_1 _14425_ (.A1(_06911_),
    .A2(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .B1(_07201_),
    .B2(_07202_),
    .C1(_01456_),
    .X(_00986_));
 sky130_fd_sc_hd__nand2_1 _14426_ (.A(_07059_),
    .B(net451),
    .Y(_07203_));
 sky130_fd_sc_hd__o21a_1 _14427_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .A2(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .B1(_07157_),
    .X(_07204_));
 sky130_fd_sc_hd__and3_1 _14428_ (.A(_07191_),
    .B(_07192_),
    .C(_07200_),
    .X(_07205_));
 sky130_fd_sc_hd__and2b_1 _14429_ (.A_N(_07196_),
    .B(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__or2_1 _14430_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_07156_),
    .X(_07207_));
 sky130_fd_sc_hd__nand2_1 _14431_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .B(_07156_),
    .Y(_07208_));
 sky130_fd_sc_hd__and2_1 _14432_ (.A(_07207_),
    .B(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__o21ai_1 _14433_ (.A1(_07204_),
    .A2(_07206_),
    .B1(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__o31a_1 _14434_ (.A1(_07209_),
    .A2(_07204_),
    .A3(_07206_),
    .B1(_01861_),
    .X(_07211_));
 sky130_fd_sc_hd__nand2_1 _14435_ (.A(_07210_),
    .B(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__a21boi_1 _14436_ (.A1(_07203_),
    .A2(_07212_),
    .B1_N(_01766_),
    .Y(_00987_));
 sky130_fd_sc_hd__xor2_1 _14437_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .B(_07156_),
    .X(_07213_));
 sky130_fd_sc_hd__a21oi_1 _14438_ (.A1(_07208_),
    .A2(_07210_),
    .B1(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__a31o_1 _14439_ (.A1(_07208_),
    .A2(_07210_),
    .A3(_07213_),
    .B1(_06926_),
    .X(_07215_));
 sky130_fd_sc_hd__o221a_1 _14440_ (.A1(_06911_),
    .A2(net518),
    .B1(_07214_),
    .B2(_07215_),
    .C1(_01456_),
    .X(_00988_));
 sky130_fd_sc_hd__xor2_1 _14441_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .B(_07157_),
    .X(_07216_));
 sky130_fd_sc_hd__and3_1 _14442_ (.A(_07209_),
    .B(_07205_),
    .C(_07213_),
    .X(_07217_));
 sky130_fd_sc_hd__and3_1 _14443_ (.A(_07172_),
    .B(_07194_),
    .C(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__a2111o_1 _14444_ (.A1(_07018_),
    .A2(_07157_),
    .B1(_07195_),
    .C1(_07204_),
    .D1(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__xor2_1 _14445_ (.A(_07216_),
    .B(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__mux2_1 _14446_ (.A0(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A1(_07220_),
    .S(_01861_),
    .X(_07221_));
 sky130_fd_sc_hd__and2_1 _14447_ (.A(_01253_),
    .B(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__clkbuf_1 _14448_ (.A(_07222_),
    .X(_00989_));
 sky130_fd_sc_hd__a22o_1 _14449_ (.A1(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ),
    .A2(_07157_),
    .B1(_07216_),
    .B2(_07219_),
    .X(_07223_));
 sky130_fd_sc_hd__xnor2_1 _14450_ (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_07157_),
    .Y(_07224_));
 sky130_fd_sc_hd__xnor2_1 _14451_ (.A(_07223_),
    .B(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__or2_1 _14452_ (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .B(_06909_),
    .X(_07226_));
 sky130_fd_sc_hd__o211a_1 _14453_ (.A1(_07059_),
    .A2(_07225_),
    .B1(_07226_),
    .C1(_01475_),
    .X(_00990_));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00000_),
    .Q(\r_i_alpha1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00001_),
    .Q(\r_i_alpha1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00002_),
    .Q(\r_i_alpha1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00003_),
    .Q(\r_i_alpha1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00004_),
    .Q(\r_i_alpha1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00005_),
    .Q(\r_i_alpha1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00006_),
    .Q(\r_i_alpha1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00007_),
    .Q(\r_i_alpha1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00008_),
    .Q(\r_i_alpha1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00009_),
    .Q(\r_i_alpha1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00010_),
    .Q(\r_i_alpha1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00011_),
    .Q(\r_i_alpha1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00012_),
    .Q(\r_i_alpha1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00013_),
    .Q(\r_i_alpha1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00014_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00015_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00016_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00017_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00018_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00019_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00020_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00021_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00022_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00023_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00024_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00025_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00026_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00027_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00028_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00029_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00030_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00031_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00032_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00033_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00034_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00035_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00036_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00037_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00038_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00039_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00040_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00041_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00042_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00043_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00044_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00045_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00046_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00047_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00048_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00049_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00050_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00051_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00052_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00053_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00054_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00055_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00056_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00057_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00058_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00059_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00060_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00061_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00062_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00063_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00064_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00065_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00066_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00067_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_2 _14522_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00068_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00069_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_in ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00070_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.i_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00071_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.i_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00072_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00073_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00074_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00075_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00076_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00077_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00078_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00079_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00080_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00081_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00082_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00083_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00084_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00085_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14540_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00086_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00087_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00088_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14543_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00089_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00090_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00091_),
    .Q(\diff1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00092_),
    .Q(\diff1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00093_),
    .Q(\diff1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00094_),
    .Q(\diff1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00095_),
    .Q(\diff1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00096_),
    .Q(\diff1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00097_),
    .Q(\diff1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00098_),
    .Q(\diff1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00099_),
    .Q(\diff1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00100_),
    .Q(\diff1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00101_),
    .Q(\diff1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00102_),
    .Q(\diff1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00103_),
    .Q(\diff1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00104_),
    .Q(\diff1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00105_),
    .Q(\diff2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00106_),
    .Q(\diff2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00107_),
    .Q(\diff2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00108_),
    .Q(\diff2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00109_),
    .Q(\diff2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00110_),
    .Q(\diff2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00111_),
    .Q(\diff2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00112_),
    .Q(\diff2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00113_),
    .Q(\diff2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00114_),
    .Q(\diff2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00115_),
    .Q(\diff2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00116_),
    .Q(\diff2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00117_),
    .Q(\diff2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00118_),
    .Q(\diff2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14573_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00119_),
    .Q(\diff2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_39_i_clk),
    .D(net2),
    .Q(diff_valid));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00120_),
    .Q(\diff1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00121_),
    .Q(\diff1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00122_),
    .Q(\diff1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00123_),
    .Q(\diff1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00124_),
    .Q(\diff3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00125_),
    .Q(\diff3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00126_),
    .Q(\diff3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00127_),
    .Q(\diff3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00128_),
    .Q(\diff3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00129_),
    .Q(\diff3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00130_),
    .Q(\diff3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00131_),
    .Q(\diff3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00132_),
    .Q(\diff3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00133_),
    .Q(\diff3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00134_),
    .Q(\diff3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00135_),
    .Q(\diff3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00136_),
    .Q(\diff3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00137_),
    .Q(\diff3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00138_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00139_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00140_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00141_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14597_ (.CLK(clknet_leaf_44_i_clk),
    .D(net402),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14598_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00143_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00144_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00145_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14601_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00146_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00147_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00148_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00149_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00150_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00151_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14607_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00152_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14608_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00153_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00154_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00155_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00156_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00157_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14613_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00158_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14614_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00159_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14615_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00160_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14616_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00161_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00162_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_4 _14618_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00163_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14619_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00164_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14620_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00165_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00166_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14622_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00167_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00168_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14624_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00169_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00170_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14626_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00171_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14627_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00172_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14628_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00173_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14629_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00174_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14630_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00175_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14631_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00176_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14632_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00177_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00178_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00179_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14635_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00180_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14636_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00181_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14637_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00182_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00183_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14639_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00184_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00185_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14641_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00186_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14642_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00187_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14643_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00188_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00189_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14645_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00190_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14646_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00191_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14647_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00192_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00193_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00194_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_50_i_clk),
    .D(net160),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00196_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00197_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_49_i_clk),
    .D(net308),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00199_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14655_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00200_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00201_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14657_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00202_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00203_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00204_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00205_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00206_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00207_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00208_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00209_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00210_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00211_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00212_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00213_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00214_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00215_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14671_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00216_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14672_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00217_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14673_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00218_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14674_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00219_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00220_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00221_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14677_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00222_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00223_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14679_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00224_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14680_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00225_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14681_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00226_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00227_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14683_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00228_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14684_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00229_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00230_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00231_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00232_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00233_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00234_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00235_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00236_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00237_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14693_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00238_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14694_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00239_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14695_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00240_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14696_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00241_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00242_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14698_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00243_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14699_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00244_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14700_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00245_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00246_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14702_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00247_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00248_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00249_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14705_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00250_),
    .Q(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_50_i_clk),
    .D(net156),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_51_i_clk),
    .D(net192),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00253_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_51_i_clk),
    .D(net301),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00255_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00256_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00257_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_50_i_clk),
    .D(net470),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00259_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00260_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00261_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14717_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00262_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14718_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00263_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00264_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_53_i_clk),
    .D(net448),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00266_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14722_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00267_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00268_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00269_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_4 _14725_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00270_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00271_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00272_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00273_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14729_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00274_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14730_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00275_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14731_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00276_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14732_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00277_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14733_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00278_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00279_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14735_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00280_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00281_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14737_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00282_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14738_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00283_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00284_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14740_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00285_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14741_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00286_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14742_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00287_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00288_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00289_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00290_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00291_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00292_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14748_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00293_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14749_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00294_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00295_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14751_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00296_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14752_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00297_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14753_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00298_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14754_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00299_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14755_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00300_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14756_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00301_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14757_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00302_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14758_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00303_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14759_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00304_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14760_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00305_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00306_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_4 _14762_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00307_),
    .Q(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00308_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_51_i_clk),
    .D(net211),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00310_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00311_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00312_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00313_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00314_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00315_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00316_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00317_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00318_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00319_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14775_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00320_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00321_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00322_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00323_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00324_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_76_i_clk),
    .D(net268),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00326_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14782_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00327_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00328_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00329_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00330_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00331_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14787_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00332_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14788_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00333_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14789_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00334_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00335_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14791_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00336_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14792_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00337_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14793_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00338_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14794_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00339_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00340_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14796_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00341_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14797_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00342_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14798_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00343_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00344_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00345_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00346_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14802_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00347_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00348_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00349_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00350_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14806_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00351_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00352_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00353_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14809_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00354_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14810_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00355_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00356_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14812_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00357_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00358_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14814_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00359_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14815_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00360_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00361_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14817_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00362_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00363_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14819_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00364_),
    .Q(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_110_i_clk),
    .D(net146),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00366_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00367_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00368_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00369_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00370_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00371_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00372_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00373_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00374_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00375_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.CLK(clknet_leaf_77_i_clk),
    .D(net604),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_77_i_clk),
    .D(net488),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00378_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00379_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14835_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00380_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00381_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00382_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00383_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14839_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00384_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00385_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00386_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00387_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00388_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00389_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14845_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00390_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14846_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00391_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14847_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00392_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00393_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00394_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14850_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00395_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14851_ (.CLK(clknet_4_7_0_i_clk),
    .D(_00396_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_4_6_0_i_clk),
    .D(_00397_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14853_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00398_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14854_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00399_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14855_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00400_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00401_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00402_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00403_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00404_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00405_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00406_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00407_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14863_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00408_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14864_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00409_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14865_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00410_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14866_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00411_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14867_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00412_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00413_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14869_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00414_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14870_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00415_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14871_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00416_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14872_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00417_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00418_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14874_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00419_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00420_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_4 _14876_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00421_),
    .Q(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_110_i_clk),
    .D(net217),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_110_i_clk),
    .D(net133),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_110_i_clk),
    .D(net142),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_110_i_clk),
    .D(net137),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_110_i_clk),
    .D(net131),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00427_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00428_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_110_i_clk),
    .D(net127),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_110_i_clk),
    .D(net125),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00431_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00432_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_109_i_clk),
    .D(net378),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00434_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00435_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00436_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00437_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00438_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00439_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00440_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14896_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00441_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00442_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00443_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00444_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00445_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00446_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00447_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14903_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00448_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14904_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00449_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00450_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00451_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14907_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00452_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00453_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14909_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00454_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14910_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00455_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00456_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00457_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14913_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00458_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00459_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00460_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00461_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00462_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00463_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00464_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00465_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14921_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00466_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14922_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00467_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14923_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00468_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00469_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14925_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00470_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14926_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00471_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14927_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00472_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00473_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14929_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00474_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14930_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00475_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00476_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00477_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00478_),
    .Q(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00479_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_110_i_clk),
    .D(net241),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00481_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00482_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_109_i_clk),
    .D(net187),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00484_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_110_i_clk),
    .D(net235),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.CLK(clknet_leaf_109_i_clk),
    .D(net180),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.CLK(clknet_leaf_109_i_clk),
    .D(net173),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00488_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.CLK(clknet_leaf_107_i_clk),
    .D(net259),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00490_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00491_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00492_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00493_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14949_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00494_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00495_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00496_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00497_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00498_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00499_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00500_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00501_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00502_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00503_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00504_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00505_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14961_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00506_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14962_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00507_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14963_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00508_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14964_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00509_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_4 _14965_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00510_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14966_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00511_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14967_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00512_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14968_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00513_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14969_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00514_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14970_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00515_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00516_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00517_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00518_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00519_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00520_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14976_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00521_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_2 _14977_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00522_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00523_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14979_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00524_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14980_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00525_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14981_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00526_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14982_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00527_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14983_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00528_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14984_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00529_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14985_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00530_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14986_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00531_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14987_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00532_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14988_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00533_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14989_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00534_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_4 _14990_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00535_),
    .Q(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00536_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00537_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00538_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00539_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00540_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00541_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00542_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00543_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00544_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_107_i_clk),
    .D(net286),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00546_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00547_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00548_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_103_i_clk),
    .D(net461),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_103_i_clk),
    .D(net464),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15006_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00551_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00552_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00553_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00554_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15010_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00555_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00556_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00557_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00558_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_4_5_0_i_clk),
    .D(_00559_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00560_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00561_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00562_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00563_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15019_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00564_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15020_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00565_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15021_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00566_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00567_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15023_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00568_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15024_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00569_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15025_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00570_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00571_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15027_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00572_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15028_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00573_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15029_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00574_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15030_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00575_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15031_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00576_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15032_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00577_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00578_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15034_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00579_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00580_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00581_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00582_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15038_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00583_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15039_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00584_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15040_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00585_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15041_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00586_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15042_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00587_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15043_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00588_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00589_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15045_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00590_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15046_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00591_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15047_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00592_),
    .Q(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15048_ (.CLK(clknet_leaf_112_i_clk),
    .D(net144),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15049_ (.CLK(clknet_leaf_111_i_clk),
    .D(net129),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15050_ (.CLK(clknet_leaf_110_i_clk),
    .D(net123),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15051_ (.CLK(clknet_leaf_111_i_clk),
    .D(net152),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15052_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00597_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15053_ (.CLK(clknet_leaf_112_i_clk),
    .D(net135),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15054_ (.CLK(clknet_leaf_112_i_clk),
    .D(net139),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15055_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00600_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15056_ (.CLK(clknet_leaf_112_i_clk),
    .D(net275),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15057_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00602_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15058_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00603_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15059_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00604_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15060_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00605_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15061_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00606_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15062_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00607_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15063_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00608_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15064_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00609_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15065_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00610_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15066_ (.CLK(clknet_leaf_117_i_clk),
    .D(net523),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_4 _15067_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00612_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15068_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00613_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15069_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00614_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15070_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00615_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15071_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00616_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15072_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00617_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15073_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00618_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15074_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00619_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00620_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00621_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15077_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00622_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15078_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00623_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15079_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00624_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15080_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00625_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15081_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00626_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15082_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00627_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15083_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00628_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15084_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00629_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15085_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00630_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00631_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00632_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00633_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00634_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00635_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00636_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00637_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00638_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00639_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15095_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00640_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15096_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00641_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15097_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00642_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_4 _15098_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00643_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15099_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00644_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15100_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00645_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15101_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00646_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00647_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00648_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00649_),
    .Q(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.CLK(clknet_leaf_111_i_clk),
    .D(net184),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.CLK(clknet_leaf_111_i_clk),
    .D(net219),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00652_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00653_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.CLK(clknet_leaf_110_i_clk),
    .D(net163),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00655_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00656_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.CLK(clknet_leaf_113_i_clk),
    .D(net343),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00658_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00659_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00660_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00661_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00662_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00663_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00664_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00665_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00666_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15122_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00667_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15123_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00668_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_4 _15124_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00669_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15125_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00670_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15126_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00671_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15127_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00672_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15128_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00673_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15129_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00674_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15130_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00675_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15131_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00676_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15132_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00677_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15133_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00678_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15134_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00679_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15135_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00680_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15136_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00681_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15137_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00682_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15138_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00683_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15139_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00684_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15140_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00685_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15141_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00686_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15142_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00687_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15143_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00688_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15144_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00689_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15145_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00690_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15146_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00691_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15147_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00692_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15148_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00693_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15149_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00694_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15150_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00695_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15151_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00696_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15152_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00697_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15153_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00698_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15154_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00699_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15155_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00700_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15156_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00701_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15157_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00702_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15158_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00703_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15159_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00704_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15160_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00705_),
    .Q(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15161_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00706_),
    .Q(\CORDIC_PE[0].genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15162_ (.CLK(clknet_leaf_111_i_clk),
    .D(net238),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15163_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00708_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15164_ (.CLK(clknet_leaf_110_i_clk),
    .D(net150),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15165_ (.CLK(clknet_leaf_110_i_clk),
    .D(net154),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15166_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00711_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15167_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00712_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15168_ (.CLK(clknet_leaf_113_i_clk),
    .D(net351),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15169_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00714_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15170_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00715_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15171_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00716_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15172_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00717_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15173_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00718_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15174_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00719_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15175_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00720_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15176_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00721_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15177_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00722_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15178_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00723_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15179_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00724_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15180_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00725_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15181_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00726_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15182_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00727_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15183_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00728_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15184_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00729_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15185_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00730_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15186_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00731_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15187_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00732_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15188_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00733_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15189_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00734_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15190_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00735_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15191_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00736_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15192_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00737_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15193_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00738_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15194_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00739_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15195_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00740_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15196_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00741_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15197_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00742_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15198_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00743_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15199_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00744_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15200_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00745_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15201_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00746_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15202_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00747_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15203_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00748_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15204_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00749_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15205_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00750_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15206_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00751_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15207_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00752_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15208_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00753_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15209_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00754_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15210_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00755_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15211_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00756_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15212_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00757_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15213_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00758_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15214_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00759_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15215_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00760_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15216_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00761_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15217_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00762_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15218_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00763_),
    .Q(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15219_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00764_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15220_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00765_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15221_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00766_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15222_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00767_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15223_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00768_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15224_ (.CLK(clknet_leaf_15_i_clk),
    .D(net436),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15225_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00770_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15226_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00771_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15227_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00772_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15228_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00773_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15229_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00774_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15230_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00775_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15231_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00776_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15232_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00777_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15233_ (.CLK(clknet_leaf_14_i_clk),
    .D(net558),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15234_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00779_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15235_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00780_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15236_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00781_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15237_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00782_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15238_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00783_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15239_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00784_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15240_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00785_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15241_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00786_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15242_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00787_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15243_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00788_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15244_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00789_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15245_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00790_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15246_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00791_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15247_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00792_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15248_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00793_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15249_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00794_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15250_ (.CLK(clknet_4_2_0_i_clk),
    .D(_00795_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15251_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00796_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15252_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00797_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15253_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00798_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15254_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00799_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15255_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00800_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15256_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00801_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15257_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00802_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15258_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00803_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15259_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00804_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15260_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00805_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15261_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00806_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15262_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00807_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15263_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00808_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15264_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00809_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15265_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00810_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15266_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00811_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15267_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00812_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15268_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00813_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15269_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00814_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15270_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00815_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15271_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00816_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15272_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00817_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15273_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00818_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15274_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00819_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15275_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00820_),
    .Q(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15276_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00821_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15277_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00822_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15278_ (.CLK(clknet_leaf_51_i_clk),
    .D(net296),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15279_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00824_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15280_ (.CLK(clknet_leaf_51_i_clk),
    .D(net457),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15281_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00826_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15282_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00827_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15283_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00828_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15284_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00829_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15285_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00830_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15286_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00831_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15287_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00832_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15288_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00833_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15289_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00834_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15290_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00835_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15291_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00836_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15292_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00837_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15293_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00838_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15294_ (.CLK(clknet_leaf_17_i_clk),
    .D(net468),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15295_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00840_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15296_ (.CLK(clknet_leaf_14_i_clk),
    .D(net612),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15297_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00842_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15298_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00843_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15299_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00844_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15300_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00845_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15301_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00846_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15302_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00847_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15303_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00848_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15304_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00849_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15305_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00850_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15306_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00851_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15307_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00852_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15308_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00853_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15309_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00854_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15310_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00855_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15311_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00856_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15312_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00857_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15313_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00858_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15314_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00859_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15315_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00860_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15316_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00861_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15317_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00862_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15318_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00863_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15319_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00864_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15320_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00865_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15321_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00866_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15322_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00867_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15323_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00868_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15324_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00869_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15325_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00870_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15326_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00871_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15327_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00872_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15328_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00873_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15329_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00874_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15330_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00875_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15331_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00876_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15332_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00877_),
    .Q(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15333_ (.CLK(clknet_leaf_23_i_clk),
    .D(net213),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15334_ (.CLK(clknet_leaf_23_i_clk),
    .D(net221),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15335_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00880_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15336_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00881_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15337_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00882_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15338_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00883_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15339_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00884_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15340_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00885_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15341_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00886_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15342_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00887_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15343_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00888_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15344_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00889_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15345_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00890_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15346_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00891_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15347_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00892_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15348_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00893_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15349_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00894_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15350_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00895_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15351_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00896_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15352_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00897_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15353_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00898_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15354_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00899_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15355_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00900_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15356_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00901_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15357_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00902_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15358_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00903_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00904_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15360_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00905_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15361_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00906_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15362_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00907_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15363_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00908_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15364_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00909_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15365_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00910_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15366_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00911_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15367_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00912_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15368_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00913_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15369_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00914_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00915_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00916_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00917_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00918_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00919_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15375_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00920_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00921_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00922_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15378_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00923_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15379_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00924_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15380_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00925_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15381_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00926_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15382_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00927_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15383_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00928_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15384_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00929_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15385_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00930_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15386_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00931_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15387_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00932_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15388_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00933_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15389_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00934_),
    .Q(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.valid_out ));
 sky130_fd_sc_hd__dfxtp_1 _15390_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00935_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15391_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00936_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15392_ (.CLK(clknet_leaf_27_i_clk),
    .D(net246),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15393_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00938_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15394_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00939_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15395_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00940_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15396_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00941_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15397_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00942_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15398_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00943_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15399_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00944_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15400_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00945_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15401_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00946_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15402_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00947_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15403_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00948_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15404_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00949_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15405_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00950_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15406_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00951_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15407_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00952_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15408_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00953_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15409_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00954_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15410_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00955_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15411_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00956_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15412_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00957_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15413_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00958_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15414_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00959_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15415_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00960_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15416_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00961_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15417_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00962_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15418_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00963_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15419_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00964_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15420_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00965_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15421_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00966_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15422_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00967_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15423_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00968_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15424_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00969_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15425_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00970_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15426_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00971_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15427_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00972_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15428_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00973_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15429_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00974_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15430_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00975_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15431_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00976_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15432_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00977_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15433_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00978_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15434_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00979_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15435_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00980_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15436_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00981_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15437_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00982_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15438_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00983_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15439_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00984_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15440_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00985_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15441_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00986_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15442_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00987_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15443_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00988_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15444_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00989_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15445_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00990_),
    .Q(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[17] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_100_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_101_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_102_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_103_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_104_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_105_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_106_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_107_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_108_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_109_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_110_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_111_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_112_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_113_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_114_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_115_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_116_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_117_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_118_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_119_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_120_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_121_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_122_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_123_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_124_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_125_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00429_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_00422_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00651_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_00879_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\diff2[6] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\diff1[9] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\diff1[5] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net83),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net96),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net80),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\diff3[5] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net110),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_00485_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00594_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_00707_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\diff2[10] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_00480_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.i_quadrant[1] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net103),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00937_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\diff3[6] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\diff3[9] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net99),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[0] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net251));
 sky130_fd_sc_hd__buf_1 hold135 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net77),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net78),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00426_),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_00489_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\diff2[15] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_00325_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_00601_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00423_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net108),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net107),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_00545_),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net291));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold175 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[1] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_00823_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_00598_),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net297));
 sky130_fd_sc_hd__buf_1 hold181 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_00254_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net92),
    .X(net302));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold186 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_01233_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net102),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_00198_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[8] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00425_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net317));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold201 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_01231_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\diff1[8] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net91),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\r_i_alpha1[9] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\r_i_alpha1[5] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net89),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[12] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_00599_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\diff1[11] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\r_i_alpha1[11] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\diff1[12] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\r_i_alpha1[7] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_00657_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\r_i_alpha1[10] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\diff1[13] ),
    .X(net345));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold229 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\diff1[6] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_01238_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_00713_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\r_i_alpha1[6] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\r_i_alpha1[13] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\diff1[1] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\diff3[16] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\diff1[15] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\r_i_alpha1[14] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\r_i_alpha1[4] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net61),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_00424_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\r_i_alpha1[12] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\r_i_alpha1[8] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net93),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net104),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net58),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net59),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net70),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net88),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net60),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\r_i_alpha1[16] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_00433_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\diff2[7] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\diff1[2] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net75),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\diff3[11] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\diff3[12] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(net74),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net94),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\r_i_alpha1[15] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_00593_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\diff3[8] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\diff1[16] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\diff2[12] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\diff3[15] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\diff2[3] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.in_alpha[2] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_00142_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\diff1[3] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_00365_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(net62),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[10] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[14] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[17] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_01248_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(net63),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(net84),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net71),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\diff2[13] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(net68),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\diff3[7] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\diff3[14] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(net64),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_01247_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net72),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_00769_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\diff2[16] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(net85),
    .X(net439));
 sky130_fd_sc_hd__buf_1 hold323 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net441));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold325 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\diff2[4] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[15] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_00709_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_00265_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net449));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold333 (.A(\diff1[0] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net90),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[16] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_00825_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[9] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[2] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_00549_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(net462));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold346 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_00550_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\diff1[17] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_00596_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_00839_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_00258_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\diff2[14] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[10] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(net81),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[0] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net480));
 sky130_fd_sc_hd__buf_1 hold364 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_00710_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_00377_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[14] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_03214_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\diff3[17] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(net79),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_00251_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[6] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[7] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[10] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net515));
 sky130_fd_sc_hd__buf_1 hold399 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_00611_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net530));
 sky130_fd_sc_hd__buf_1 hold414 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[13] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[4] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[10] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_00195_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[14] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[0] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_00778_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[12] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[11] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[7] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_00654_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_x[9] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[6] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[15] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[7] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[13] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[7] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[14] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[9] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_00376_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_x[15] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[15] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(net87),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_06297_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_00841_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[3] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\CORDIC_PE[7].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net86),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[5] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_x[1] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_x[11] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[10] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_x[5] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_x[17] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net106),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[13] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[12] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_x[3] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[11] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_y[1] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[8] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\CORDIC_PE[3].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_alpha[8] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_y[4] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\CORDIC_PE[13].genblk1.genblk1.cordic_engine_inst.out_y[4] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_y[8] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_x[4] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[17] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\CORDIC_PE[9].genblk1.genblk1.cordic_engine_inst.out_alpha[11] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_y[13] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\CORDIC_PE[11].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net98),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_y[0] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[16] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net105),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_00487_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00595_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net100),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\r_i_alpha1[17] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_00486_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\diff1[10] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net95),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_00650_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net109),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\CORDIC_PE[5].genblk1.genblk1.cordic_engine_inst.out_alpha[2] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_00483_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\diff1[14] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\diff3[4] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\diff1[7] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\CORDIC_PE[1].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00252_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net101),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\diff2[11] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\diff2[9] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\diff2[5] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00430_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net97),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\diff3[10] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\diff2[8] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\diff3[13] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[4] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\diff1[4] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_alpha[0] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[3] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\CORDIC_PE[0].genblk1.cordic_engine_inst.i_quadrant[0] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_alpha[5] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\CORDIC_PE[10].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net111),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_alpha[1] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\CORDIC_PE[2].genblk1.genblk1.cordic_engine_inst.out_quadrant[1] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00309_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\CORDIC_PE[12].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_00878_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net82),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\CORDIC_PE[14].genblk1.genblk1.cordic_engine_inst.out_alpha[6] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\CORDIC_PE[4].genblk1.genblk1.cordic_engine_inst.out_quadrant[0] ),
    .X(net216));
 sky130_fd_sc_hd__buf_1 input1 (.A(i_rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(in_alpha[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(in_alpha[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in_alpha[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(in_alpha[2]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(in_alpha[3]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(in_alpha[4]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(in_alpha[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(in_alpha[6]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(in_alpha[7]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(in_alpha[8]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(i_valid_in),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(in_alpha[9]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(in_x[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in_x[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in_x[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in_x[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(in_x[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in_x[14]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(in_x[15]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(in_x[16]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(in_x[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(in_alpha[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(in_x[1]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in_x[2]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(in_x[3]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(in_x[4]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(in_x[5]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(in_x[6]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(in_x[7]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(in_x[8]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in_x[9]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(in_y[0]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(in_alpha[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in_y[10]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in_y[11]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in_y[12]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(in_y[13]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(in_y[14]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(in_y[15]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(in_y[16]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(in_y[17]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(in_y[1]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(in_y[2]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(in_alpha[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(in_y[3]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in_y[4]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(in_y[5]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(in_y[6]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in_y[7]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(in_y[8]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in_y[9]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input6 (.A(in_alpha[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(in_alpha[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(in_alpha[14]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(in_alpha[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 max_cap114 (.A(_05015_),
    .X(net114));
 sky130_fd_sc_hd__buf_1 max_cap117 (.A(_03700_),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(out_sintheta[15]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(out_sintheta[16]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(out_sintheta[17]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(out_sintheta[1]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(out_sintheta[2]));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(out_sintheta[3]));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(out_sintheta[4]));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(out_sintheta[5]));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(out_sintheta[6]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(out_sintheta[7]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(out_sintheta[8]));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(out_sintheta[9]));
 sky130_fd_sc_hd__clkbuf_4 output57 (.A(net57),
    .X(o_valid_out));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(out_alpha[0]));
 sky130_fd_sc_hd__clkbuf_4 output59 (.A(net59),
    .X(out_alpha[10]));
 sky130_fd_sc_hd__clkbuf_4 output60 (.A(net60),
    .X(out_alpha[11]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(out_alpha[12]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(out_alpha[13]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(out_alpha[14]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(out_alpha[15]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(out_alpha[16]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(out_alpha[17]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(out_alpha[1]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(out_alpha[2]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(out_alpha[3]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(out_alpha[4]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(out_alpha[5]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(out_alpha[6]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(out_alpha[7]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(out_alpha[8]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(out_alpha[9]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(out_costheta[0]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(out_costheta[10]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(out_costheta[11]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(out_costheta[12]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(out_costheta[13]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(out_costheta[14]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(out_costheta[15]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(out_costheta[16]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(out_costheta[17]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(out_costheta[1]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(out_costheta[2]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(out_costheta[3]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(out_costheta[4]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(out_costheta[5]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(out_costheta[6]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(out_costheta[7]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(out_costheta[8]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(out_costheta[9]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(out_sintheta[0]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .X(out_sintheta[10]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(out_sintheta[11]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(out_sintheta[12]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(out_sintheta[13]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(out_sintheta[14]));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(\CORDIC_PE[6].genblk1.genblk1.cordic_engine_inst.out_y[9] ),
    .X(net120));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(_05236_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_04632_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(\CORDIC_PE[8].genblk1.genblk1.cordic_engine_inst.out_x[12] ),
    .X(net653));
 sky130_fd_sc_hd__buf_1 wire113 (.A(_06051_),
    .X(net113));
 sky130_fd_sc_hd__buf_1 wire115 (.A(_04269_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 wire116 (.A(_06805_),
    .X(net116));
endmodule

