* NGSPICE file created from cordic_tt_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

.subckt cordic_tt_top VGND VPWR i_clk i_rst_n i_valid_in in_alpha[0] in_alpha[10]
+ in_alpha[11] in_alpha[12] in_alpha[13] in_alpha[14] in_alpha[15] in_alpha[16] in_alpha[17]
+ in_alpha[1] in_alpha[2] in_alpha[3] in_alpha[4] in_alpha[5] in_alpha[6] in_alpha[7]
+ in_alpha[8] in_alpha[9] in_x[0] in_x[10] in_x[11] in_x[12] in_x[13] in_x[14] in_x[15]
+ in_x[16] in_x[17] in_x[1] in_x[2] in_x[3] in_x[4] in_x[5] in_x[6] in_x[7] in_x[8]
+ in_x[9] in_y[0] in_y[10] in_y[11] in_y[12] in_y[13] in_y[14] in_y[15] in_y[16] in_y[17]
+ in_y[1] in_y[2] in_y[3] in_y[4] in_y[5] in_y[6] in_y[7] in_y[8] in_y[9] o_valid_out
+ out_alpha[0] out_alpha[10] out_alpha[11] out_alpha[12] out_alpha[13] out_alpha[14]
+ out_alpha[15] out_alpha[16] out_alpha[17] out_alpha[1] out_alpha[2] out_alpha[3]
+ out_alpha[4] out_alpha[5] out_alpha[6] out_alpha[7] out_alpha[8] out_alpha[9] out_costheta[0]
+ out_costheta[10] out_costheta[11] out_costheta[12] out_costheta[13] out_costheta[14]
+ out_costheta[15] out_costheta[16] out_costheta[17] out_costheta[1] out_costheta[2]
+ out_costheta[3] out_costheta[4] out_costheta[5] out_costheta[6] out_costheta[7]
+ out_costheta[8] out_costheta[9] out_sintheta[0] out_sintheta[10] out_sintheta[11]
+ out_sintheta[12] out_sintheta[13] out_sintheta[14] out_sintheta[15] out_sintheta[16]
+ out_sintheta[17] out_sintheta[1] out_sintheta[2] out_sintheta[3] out_sintheta[4]
+ out_sintheta[5] out_sintheta[6] out_sintheta[7] out_sintheta[8] out_sintheta[9]
XFILLER_0_94_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09671_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03080_ VGND
+ VGND VPWR VPWR _03082_ sky130_fd_sc_hd__or2_1
X_08622_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _02152_ sky130_fd_sc_hd__inv_2
X_08553_ _01867_ _02089_ _02090_ _01552_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07504_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _01122_ _01156_
+ _01046_ _01072_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__a221o_1
X_08484_ _02025_ _02026_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07435_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _01159_ _01164_
+ _01168_ _01059_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__o221a_1
XFILLER_0_92_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07366_ _01105_ _01106_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09105_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__and2b_1
X_07297_ _01015_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_4
X_09036_ _02513_ _02508_ _02516_ _02369_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold340 _00825_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold351 _00839_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold362 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold373 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ _03313_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__clkbuf_1
X_09869_ _03237_ net532 _03251_ _03254_ _03013_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11900_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _05027_ VGND
+ VGND VPWR VPWR _05028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12880_ _05853_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__clkbuf_4
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04930_ VGND
+ VGND VPWR VPWR _04966_ sky130_fd_sc_hd__or2_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ clknet_leaf_35_i_clk _00096_ VGND VGND VPWR VPWR diff1\[9\] sky130_fd_sc_hd__dfxtp_1
X_11762_ _04795_ _04904_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nand2_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13501_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06407_
+ _06408_ _06285_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__o221a_1
X_10713_ net157 _03997_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__or2_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14481_ clknet_leaf_25_i_clk _00027_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04841_ VGND
+ VGND VPWR VPWR _04842_ sky130_fd_sc_hd__xnor2_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13432_ _06069_ _06348_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10644_ _03935_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10575_ _03860_ _03867_ _03865_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__o21a_1
X_13363_ _06286_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15102_ clknet_leaf_118_i_clk _00647_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12314_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05384_ VGND
+ VGND VPWR VPWR _05385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13294_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _06218_
+ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15033_ clknet_leaf_97_i_clk _00578_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12245_ _05290_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12176_ _05262_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _05263_ sky130_fd_sc_hd__and2_4
X_11127_ _04349_ _04353_ _04357_ _04047_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_120_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_120_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11058_ _04295_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10009_ _03364_ _03374_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__o21ai_1
X_14817_ clknet_leaf_74_i_clk _00362_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_149_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14748_ clknet_leaf_72_i_clk _00293_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_80_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14679_ clknet_leaf_63_i_clk _00224_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_74_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07984_ _01539_ net613 _01583_ _01586_ _01513_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__o221a_1
X_09723_ _02748_ _03128_ _03129_ _03058_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__o211a_1
X_09654_ _02844_ net573 _03065_ _03066_ _03013_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08605_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[0\]
+ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nor2_1
X_09585_ _02962_ _03002_ _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__a21bo_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _02059_ _02067_ _02073_ _01924_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\] _02010_ VGND VGND VPWR
+ VPWR _02011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07418_ _01019_ _01152_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__nor2_1
X_08398_ _01877_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07349_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _01082_ VGND
+ VGND VPWR VPWR _01092_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10360_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _03680_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09019_ _02501_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10291_ _03606_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__clkbuf_4
X_12030_ _01250_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net298 sky130_fd_sc_hd__buf_1
Xhold192 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR VPWR
+ net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13981_ _06815_ _06817_ _06814_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_52_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12932_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05905_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__nand2_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ clknet_leaf_45_i_clk _00147_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11814_ _04755_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] VGND
+ VGND VPWR VPWR _04951_ sky130_fd_sc_hd__and2_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _05800_ _05801_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__and2_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ clknet_leaf_39_i_clk _00079_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11745_ _04888_ _04882_ _04883_ _04757_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__o31a_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14464_ clknet_leaf_36_i_clk _00010_ VGND VGND VPWR VPWR r_i_alpha1\[14\] sky130_fd_sc_hd__dfxtp_1
X_11676_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _04824_
+ _04823_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06332_ VGND
+ VGND VPWR VPWR _06333_ sky130_fd_sc_hd__nand2_1
X_10627_ _03650_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14395_ _07175_ _07176_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13346_ _06210_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _06203_ _06273_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__o211a_1
X_10558_ _03858_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13277_ _06213_ _06214_ _05928_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__a21oi_1
X_10489_ _03789_ _03792_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__o21ba_1
X_15016_ clknet_leaf_101_i_clk _00561_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12228_ _05308_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__and2_1
X_12159_ _05246_ _05247_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09370_ _02812_ _02813_ _02409_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08321_ _01867_ _01884_ _01885_ _01552_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08252_ _01680_ _01662_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08183_ _01556_ _01771_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07967_ _01554_ _01569_ _01570_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__a21o_1
X_09706_ _03101_ _03112_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__a21o_1
X_07898_ _01252_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__buf_6
X_09637_ _03047_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09568_ _02988_ _02981_ _02983_ _02745_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08519_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[10\] _02058_ VGND VGND VPWR
+ VPWR _02059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09499_ _02907_ _02901_ _02914_ _02925_ _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a32o_1
X_11530_ _04708_ _04700_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11461_ _04442_ _04644_ _04645_ _04456_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13200_ _06150_ _06146_ _06147_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__o31a_1
X_10412_ _03724_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11392_ _04585_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__clkbuf_1
X_14180_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _06984_ _06934_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13131_ _05841_ _06088_ _06089_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__or3_1
X_10343_ net537 _03665_ _03606_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13062_ _06025_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__xor2_1
X_10274_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] _03609_
+ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12013_ _05127_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
X_13964_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] net116 _06807_
+ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__a21o_1
X_12915_ _05566_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _05890_ _05900_
+ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__o41a_1
XFILLER_0_88_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13895_ _06556_ _06745_ _06746_ _06747_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12846_ net148 _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__or2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05781_ VGND
+ VGND VPWR VPWR _05787_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ clknet_leaf_33_i_clk _00062_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
X_11728_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04873_ VGND
+ VGND VPWR VPWR _04874_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14447_ _01253_ _07221_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11659_ _04445_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04807_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__o31a_1
XFILLER_0_142_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14378_ _07161_ _07155_ _07158_ _01861_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13329_ _05927_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _06247_ _06258_
+ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__o41a_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08870_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _02363_
+ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__or2_1
X_07821_ net9 _01445_ net10 VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__o21ai_1
X_07752_ _01399_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__nand2_1
X_07683_ net326 _01351_ _01000_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09422_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _02856_ VGND
+ VGND VPWR VPWR _02857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09353_ _02754_ net395 _02749_ _02799_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08304_ _01867_ net159 _01823_ _01872_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09284_ _02740_ _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08235_ _01672_ _01814_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08166_ _01750_ _01738_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08097_ _01689_ _01690_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__nor2_4
XFILLER_0_113_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08999_ _02342_ _02483_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10961_ _04208_ _04209_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ _03993_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__a2bb2o_1
X_12700_ _05703_ _05708_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__a21o_1
X_13680_ _06562_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__clkbuf_4
X_10892_ _04145_ _04146_ _03997_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12631_ _05653_ _05654_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_54_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15350_ clknet_leaf_48_i_clk _00895_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_12562_ _05290_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14301_ _07095_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
X_11513_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ _04671_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND
+ VPWR VPWR _04693_ sky130_fd_sc_hd__or4b_1
X_15281_ clknet_leaf_16_i_clk _00826_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12493_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05536_
+ _05489_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14232_ _07029_ _07032_ _07030_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11444_ _04237_ _04621_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14163_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06973_
+ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__or2_1
X_11375_ _04569_ _04563_ _04566_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13114_ _06071_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__xnor2_1
X_10326_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03644_
+ _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__o21ai_1
X_14094_ _06917_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__or2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _06010_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__o21ai_1
X_10257_ _03599_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10188_ _03105_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14996_ clknet_leaf_108_i_clk _00541_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13947_ _06501_ _06792_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13878_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND
+ VGND VPWR VPWR _06733_ sky130_fd_sc_hd__or2_1
X_12829_ _05808_ _05816_ _05830_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08020_ _01589_ _01591_ _01603_ _01618_ _01619_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__a311o_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09971_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03342_ VGND
+ VGND VPWR VPWR _03343_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08922_ _02387_ net449 _02412_ _02413_ _02414_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08853_ _02354_ _02355_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07804_ _01435_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__nor2_1
X_08784_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[16\] _02299_ VGND VGND VPWR
+ VPWR _02300_ sky130_fd_sc_hd__xor2_1
X_07735_ net19 _01385_ _01344_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__a21oi_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ _00992_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_4
X_09405_ _02841_ _02842_ _02843_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07597_ _01283_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09336_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR _02785_ sky130_fd_sc_hd__inv_2
X_09267_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _02117_ _02712_
+ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08218_ _01598_ _01800_ _01612_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09198_ _02662_ _02663_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08149_ _01738_ _01739_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11160_ net166 _04379_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10111_ _03467_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__and2b_1
X_11091_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04325_ _04326_
+ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__or3_1
X_10042_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03391_ _03407_
+ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__o21ai_1
Xhold30 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ clknet_leaf_84_i_clk _00395_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold63 _00486_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND VGND
+ VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 diff1\[4\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _00878_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13801_ _06658_ _06659_ _06664_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__o21ai_2
X_14781_ clknet_leaf_75_i_clk _00326_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11993_ _05102_ _05107_ _05103_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__o21ba_1
X_13732_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06600_
+ _06587_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__a21oi_2
X_10944_ _04191_ _04193_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13663_ _06543_ _06545_ _06549_ _06200_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__a31o_1
X_10875_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15402_ clknet_leaf_37_i_clk _00947_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12614_ _05636_ _05638_ _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13594_ _06489_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__nand2_1
X_15333_ clknet_leaf_23_i_clk net213 VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12545_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05578_ VGND
+ VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15264_ clknet_leaf_10_i_clk _00809_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12476_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _05516_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__or3_1
XFILLER_0_81_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14215_ _07020_ _06934_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__mux2_1
X_11427_ _04601_ _04606_ _04614_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a21o_1
X_15195_ clknet_leaf_0_i_clk _00740_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _06647_ _06960_ _06962_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__o21a_1
X_11358_ _04468_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10309_ _03630_ _03636_ _03606_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__a21o_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14077_ _01862_ _01010_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__or2_1
X_11289_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _04490_ VGND
+ VGND VPWR VPWR _04492_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _05986_ _05999_ _05994_ _05992_ _05984_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14979_ clknet_leaf_89_i_clk _00524_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_07520_ net421 net323 _01013_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__mux2_1
X_07451_ _01051_ _01033_ _01034_ _01081_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07382_ _01047_ _01119_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09121_ _02497_ _02593_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09052_ _02314_ _02531_ _02532_ _02260_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08003_ _01589_ _01593_ _01588_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold500 net86 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold511 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09954_ _03314_ _03320_ _03318_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08905_ _01959_ _02399_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__o21ba_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _02851_ _03265_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__o21a_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _02341_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__buf_2
X_08767_ _01881_ _02283_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__nand2_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ net397 _01334_ _01358_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__mux2_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[10\] _02220_ VGND VGND VPWR
+ VPWR _02221_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07649_ diff2\[16\] _01269_ _01271_ diff3\[16\] _01324_ VGND VGND VPWR VPWR _01325_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10660_ _03946_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09319_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10591_ _03888_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12330_ _05397_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12261_ _05338_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14000_ _06838_ _06834_ _06836_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__and3b_1
XFILLER_0_121_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11212_ _04391_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__nand2_1
X_12192_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05164_ _05277_
+ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__a21o_1
X_11143_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04011_ _04371_
+ _04372_ _04360_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput64 net64 VGND VGND VPWR VPWR out_alpha[15] sky130_fd_sc_hd__clkbuf_4
Xoutput75 net75 VGND VGND VPWR VPWR out_alpha[9] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR out_costheta[2] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 VGND VGND VPWR VPWR out_sintheta[12] sky130_fd_sc_hd__clkbuf_4
X_11074_ _04297_ _04305_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__nor2_1
X_14902_ clknet_leaf_83_i_clk _00447_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10025_ _03207_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__and2_1
X_14833_ clknet_leaf_76_i_clk _00378_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14764_ clknet_leaf_51_i_clk net211 VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11976_ _04770_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _05097_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13715_ _06565_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _06591_ _06592_ _06526_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__o221a_1
X_10927_ _04169_ _04174_ _04175_ _04176_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14695_ clknet_leaf_61_i_clk _00240_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13646_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06514_ VGND
+ VGND VPWR VPWR _06536_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10858_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04116_ _03996_
+ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13577_ _06472_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10789_ _04054_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__or2b_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15316_ clknet_leaf_22_i_clk _00861_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12528_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _05566_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15247_ clknet_leaf_8_i_clk _00792_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12459_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND VPWR
+ VPWR _05508_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15178_ clknet_leaf_115_i_clk _00723_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14129_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _06948_
+ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09670_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03080_ VGND
+ VGND VPWR VPWR _03081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08621_ _02145_ _02143_ _02149_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08552_ _01873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _02090_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07503_ _01022_ _01152_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__nor2_1
X_08483_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\] _02008_ _01879_ VGND
+ VGND VPWR VPWR _02026_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07434_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _01051_ _01052_
+ _01167_ _01057_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07365_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _01096_ VGND
+ VGND VPWR VPWR _01106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09104_ _02321_ net291 _02381_ _02578_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07296_ _01043_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09035_ _02513_ _02508_ _02516_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold330 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold341 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\] VGND VGND VPWR VPWR
+ net458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold385 diff3\[17\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09937_ _03312_ _03118_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__and2b_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _02851_ _03252_ _03253_ _03201_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a31o_1
X_08819_ _02326_ _02327_ _02322_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__o21ai_1
X_09799_ _02851_ _03193_ _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__and3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _04771_ net589 _04963_ _04964_ _04965_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__o221a_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04864_ _04903_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _06405_ _06406_ _06216_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__a21o_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__clkbuf_4
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ clknet_leaf_25_i_clk _00026_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11692_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _04841_ sky130_fd_sc_hd__o21ba_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13431_ _06346_ _06347_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ _06200_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10643_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03934_ VGND
+ VGND VPWR VPWR _03936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06280_
+ _06235_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a21o_1
X_10574_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03871_ VGND
+ VGND VPWR VPWR _03873_ sky130_fd_sc_hd__or2_1
X_15101_ clknet_leaf_118_i_clk _00646_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12313_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05375_ _05164_
+ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13293_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _06214_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__or3_1
X_15032_ clknet_leaf_91_i_clk _00577_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12244_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05323_ _01249_
+ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12175_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05261_ VGND
+ VGND VPWR VPWR _05262_ sky130_fd_sc_hd__xnor2_1
X_11126_ _04349_ _04353_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a21oi_1
X_11057_ _04292_ _04294_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10008_ _03375_ _03366_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__a21o_1
X_14816_ clknet_leaf_68_i_clk _00361_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11959_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05081_ VGND
+ VGND VPWR VPWR _05082_ sky130_fd_sc_hd__xor2_1
X_14747_ clknet_leaf_73_i_clk _00292_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14678_ clknet_leaf_63_i_clk _00223_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13629_ _06201_ _06520_ _06521_ _06459_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07983_ _01556_ _01585_ _01480_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09722_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND
+ VGND VPWR VPWR _03129_ sky130_fd_sc_hd__or2_1
X_09653_ _03063_ _03064_ _02747_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__a21o_1
X_08604_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[0\]
+ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__and2_1
X_09584_ _02981_ _03003_ _02994_ _02993_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08535_ _02059_ _02067_ _02073_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08466_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\] _02009_ VGND VGND VPWR
+ VPWR _02010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07417_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _01143_ VGND
+ VGND VPWR VPWR _01152_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08397_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[15\] _01949_ VGND VGND
+ VPWR VPWR _01950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07348_ _01019_ _01090_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07279_ _01019_ _01020_ _01027_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09018_ _02488_ _02494_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__nand2_1
X_10290_ _03607_ net298 _03620_ _03622_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold160 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
X_13980_ _06820_ _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__nand2_1
X_12931_ _05871_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _05913_ _05914_ _05910_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__o221a_1
X_12862_ _05854_ net435 _05847_ _05856_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__o211a_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _04771_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04949_
+ _04950_ _04788_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__o221a_1
X_14601_ clknet_leaf_46_i_clk _00146_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05781_ VGND
+ VGND VPWR VPWR _05801_ sky130_fd_sc_hd__xor2_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ clknet_leaf_39_i_clk _00078_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11744_ _04882_ _04883_ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__o21ai_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ clknet_leaf_36_i_clk _00009_ VGND VGND VPWR VPWR r_i_alpha1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11675_ _04773_ net522 _04826_ _04827_ _04788_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13414_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06324_ VGND
+ VGND VPWR VPWR _06332_ sky130_fd_sc_hd__nor2_1
X_10626_ _03862_ _03879_ _03904_ _03919_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__or4_4
X_14394_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _07157_ _07172_
+ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13345_ _06268_ _06271_ _06272_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__o21ai_1
X_10557_ _03535_ _03857_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13276_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10488_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03796_ VGND
+ VGND VPWR VPWR _03797_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15015_ clknet_leaf_100_i_clk _00560_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12227_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05291_ _05295_
+ _05292_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _05245_ VGND
+ VGND VPWR VPWR _05247_ sky130_fd_sc_hd__or2b_1
X_11109_ _04010_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _04344_ sky130_fd_sc_hd__or2_1
X_12089_ _04829_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05182_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ _01873_ net618 VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08251_ _01330_ _01698_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08182_ _01769_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07966_ net30 net48 VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__and2b_1
X_09705_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03098_ VGND
+ VGND VPWR VPWR _03113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07897_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\] _01509_ _01480_
+ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__a21o_1
X_09636_ _02924_ _03049_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__xnor2_1
X_09567_ _02981_ _02983_ _02988_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08518_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\] _02057_ VGND VGND VPWR
+ VPWR _02058_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09498_ _02924_ _02913_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08449_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[4\] _01994_ VGND VGND VPWR
+ VPWR _01995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11460_ _04444_ net493 VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10411_ _03699_ _03725_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__a21o_1
X_11391_ _04468_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13130_ _06081_ _06075_ _06087_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_61_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10342_ net526 _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__nor2_1
X_13061_ _06027_ _06028_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__and2_1
X_10273_ _03607_ net141 _03568_ _03612_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12012_ _04758_ _02310_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__and2_1
X_13963_ _06806_ _06292_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__mux2_2
X_12914_ _05567_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _05895_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__nand3_1
XFILLER_0_88_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13894_ _04455_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__clkbuf_4
X_12845_ _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__clkbuf_4
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05781_ VGND
+ VGND VPWR VPWR _05786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04864_ _04794_
+ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14515_ clknet_leaf_32_i_clk _00061_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11658_ _04445_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04808_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14446_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _07220_ _01861_
+ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10609_ _03862_ _03879_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14377_ _07155_ _07158_ _07161_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11589_ _04756_ net143 _04387_ _04759_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13328_ _05928_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _06253_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13259_ _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07820_ net9 net10 _01445_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07751_ _01003_ net7 _01395_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__or3_2
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07682_ _01349_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09421_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09352_ _02755_ _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__nand2_1
X_08303_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _01870_
+ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09283_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _02726_ VGND
+ VGND VPWR VPWR _02741_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08234_ _01638_ _01810_ _01636_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08165_ _01749_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_51_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08096_ net24 net42 VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08998_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ _02442_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__or4_2
X_07949_ _01485_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10960_ _04204_ _04207_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__nor2_1
X_09619_ _03034_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
X_10891_ _04145_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__and2_1
X_12630_ _05655_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12561_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05594_ _05489_
+ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11512_ _04691_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__buf_6
X_14300_ _01253_ _07094_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15280_ clknet_leaf_51_i_clk net457 VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12492_ _05534_ _05535_ _05526_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14231_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _07023_ VGND
+ VGND VPWR VPWR _07035_ sky130_fd_sc_hd__xnor2_1
X_11443_ _04629_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_19_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14162_ _06928_ net320 _06975_ _06976_ _06922_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11374_ _04563_ _04566_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13113_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06072_ VGND
+ VGND VPWR VPWR _06073_ sky130_fd_sc_hd__xnor2_1
X_10325_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14093_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND VPWR
+ VPWR _06918_ sky130_fd_sc_hd__a21oi_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _05842_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] VGND
+ VGND VPWR VPWR _06014_ sky130_fd_sc_hd__and2_1
X_10256_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _03572_ VGND
+ VGND VPWR VPWR _03600_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03537_ VGND
+ VGND VPWR VPWR _03538_ sky130_fd_sc_hd__xor2_2
X_14995_ clknet_leaf_109_i_clk _00540_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13946_ _06554_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _06790_
+ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__a22o_1
X_13877_ _06562_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__buf_2
X_12828_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _05789_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _05767_ _05769_ _05770_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__o21ai_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14429_ _07196_ _07205_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__and2b_1
XFILLER_0_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09970_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _03205_ _03331_
+ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08921_ _02308_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08852_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR _02356_ sky130_fd_sc_hd__inv_2
X_07803_ net4 _01431_ net5 VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__a21oi_1
X_08783_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[17\] _02296_ _02298_ VGND
+ VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07734_ net19 _01385_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__or2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07665_ _00991_ _01334_ net16 VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__o21a_1
X_09404_ _02751_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _01794_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__o21ai_1
X_07596_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[5\] _01281_ _01282_ VGND
+ VGND VPWR VPWR _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ _02409_ _02783_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09266_ _02725_ _01958_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08217_ _01597_ _01796_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09197_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _02661_ VGND
+ VGND VPWR VPWR _02663_ sky130_fd_sc_hd__or2_1
X_08148_ _01722_ _01731_ _01720_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08079_ _01647_ _01673_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__o21a_1
X_10110_ _03035_ _03466_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nand2_1
X_11090_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04205_ net115
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR VPWR
+ _04326_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_101_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10041_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR _03407_ sky130_fd_sc_hd__inv_2
Xhold20 _00425_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_quadrant\[1\] VGND VGND VPWR
+ VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 net98 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 diff1\[10\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 _00252_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _06662_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__and2_1
Xhold86 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND VPWR
+ VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 net82 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _05110_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
X_14780_ clknet_leaf_76_i_clk net268 VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10943_ _04191_ _04193_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__nor2_1
X_13731_ _06293_ _06605_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10874_ _04085_ _04092_ _04113_ _04130_ _04123_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__a2111o_1
X_13662_ _06543_ _06545_ _06549_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15401_ clknet_leaf_37_i_clk _00946_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12613_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _05641_ VGND
+ VGND VPWR VPWR _05642_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13593_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06488_ VGND
+ VGND VPWR VPWR _06490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12544_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05578_ VGND
+ VGND VPWR VPWR _05579_ sky130_fd_sc_hd__nor2_1
X_15332_ clknet_leaf_19_i_clk _00877_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12475_ _05489_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__clkbuf_4
X_15263_ clknet_leaf_10_i_clk _00808_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11426_ _04605_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _04614_ sky130_fd_sc_hd__and2b_1
X_14214_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _07018_ _06934_
+ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__o21ai_1
X_15194_ clknet_leaf_0_i_clk _00739_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14145_ _06646_ _06961_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__nand2_1
X_11357_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04554_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10308_ _03630_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__nor2_1
X_14076_ _06904_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__clkbuf_4
X_11288_ _04490_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _04491_ sky130_fd_sc_hd__and2b_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _05964_ _05971_ _05972_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__o21ai_1
X_10239_ _03584_ _03585_ _03186_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__and3b_1
X_14978_ clknet_leaf_93_i_clk _00523_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13929_ _06561_ net324 _06678_ _06776_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07450_ _01044_ net439 _01180_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07381_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _01105_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__o21ai_1
X_09120_ _02319_ _02589_ _02590_ _02592_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09051_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _02532_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08002_ _01597_ _01598_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold501 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold512 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND VPWR VPWR
+ net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND VGND VPWR
+ VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09953_ _03325_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__and2b_1
X_08904_ _01958_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _02393_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__and3_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _03253_ _03266_ _02850_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__o21ai_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _02341_ sky130_fd_sc_hd__inv_2
X_08766_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\] _02249_ VGND VGND VPWR VPWR
+ _02283_ sky130_fd_sc_hd__or4_4
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ net466 _01333_ _01375_ _01376_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__o22a_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\] _02208_ _01880_ VGND
+ VGND VPWR VPWR _02220_ sky130_fd_sc_hd__o21a_1
X_07648_ diff2\[17\] diff1\[16\] VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__and2_1
X_07579_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[3\] _01267_ _01255_ VGND
+ VGND VPWR VPWR _01268_ sky130_fd_sc_hd__mux2_1
X_09318_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _02769_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10590_ _03535_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09249_ _02333_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND
+ VGND VPWR VPWR _02710_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12260_ _05290_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11211_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _04423_
+ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__xnor2_1
X_12191_ _05163_ _05276_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__a21oi_1
X_11142_ _04364_ _04366_ _04370_ _04047_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__a31o_1
Xoutput65 net65 VGND VGND VPWR VPWR out_alpha[16] sky130_fd_sc_hd__clkbuf_4
Xoutput76 net76 VGND VGND VPWR VPWR out_costheta[0] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 VGND VGND VPWR VPWR out_costheta[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11073_ _04279_ _04274_ _04286_ _04290_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__o31ai_2
Xoutput98 net98 VGND VGND VPWR VPWR out_sintheta[13] sky130_fd_sc_hd__clkbuf_4
X_14901_ clknet_leaf_87_i_clk _00446_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10024_ _03370_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__or2_1
X_14832_ clknet_leaf_77_i_clk net488 VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14763_ clknet_leaf_51_i_clk _00308_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11975_ _05092_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13714_ _06590_ _06588_ _06589_ _06569_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__a31o_1
X_10926_ _04169_ _04174_ _04175_ _04176_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__a41o_1
X_14694_ clknet_leaf_57_i_clk _00239_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10857_ _04113_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__xor2_1
X_13645_ _06529_ _06531_ _06528_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_39_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _04041_ _04035_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__a31o_1
X_13576_ _06450_ _06473_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__o21a_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_15_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15315_ clknet_leaf_18_i_clk _00860_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12527_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05561_
+ _05560_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15246_ clknet_leaf_12_i_clk _00791_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12458_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND VPWR
+ VPWR _05507_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11409_ _04592_ _04594_ _04598_ _04396_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12389_ _05451_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15177_ clknet_leaf_114_i_clk _00722_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14128_ _06647_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _06940_ _06947_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14059_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _06845_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__o41a_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _02145_ _02143_ _02149_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__o21bai_2
X_08551_ _02082_ _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07502_ _01015_ net477 _01218_ _01219_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08482_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR VPWR
+ _02025_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07433_ _01165_ _01166_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07364_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _01096_ VGND
+ VGND VPWR VPWR _01105_ sky130_fd_sc_hd__or2_4
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09103_ _02576_ _02577_ _02322_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07295_ net370 _01042_ _01013_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09034_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _02515_ VGND
+ VGND VPWR VPWR _02516_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold320 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND VPWR
+ VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold331 _00265_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\] VGND VGND VPWR VPWR
+ net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _00258_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net481 sky130_fd_sc_hd__buf_1
Xhold375 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold397 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[10\] VGND VGND VPWR VPWR
+ net514 sky130_fd_sc_hd__dlygate4sd3_1
X_09936_ _03182_ _03309_ _03310_ _03311_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__o31a_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _03244_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__nand3_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _02324_ _02325_ _01959_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a21oi_1
X_09798_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nand2_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _02263_ _02266_ _01866_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__or4_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _03996_ sky130_fd_sc_hd__buf_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11691_ _04832_ _04836_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__nor2_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10642_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03934_ VGND
+ VGND VPWR VPWR _03935_ sky130_fd_sc_hd__and2_1
X_13430_ _06338_ _06344_ _06345_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13361_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06279_
+ _06235_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10573_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03871_ VGND
+ VGND VPWR VPWR _03872_ sky130_fd_sc_hd__nand2_2
X_15100_ clknet_leaf_118_i_clk _00645_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_12312_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR _05383_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13292_ _06223_ net516 _06226_ _06227_ _06197_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15031_ clknet_leaf_91_i_clk _00576_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12243_ _05319_ _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12174_ _05260_ _05163_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__and2_4
X_11125_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04338_ VGND
+ VGND VPWR VPWR _04357_ sky130_fd_sc_hd__xor2_2
X_11056_ _04292_ _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10007_ _03375_ _03366_ _03359_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14815_ clknet_leaf_70_i_clk _00360_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14746_ clknet_leaf_73_i_clk _00291_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11958_ _05072_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10909_ _04155_ _04159_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__or2b_1
XFILLER_0_157_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14677_ clknet_leaf_63_i_clk _00222_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_11889_ _05014_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13628_ _06204_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _06521_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13559_ _06201_ _06457_ _06458_ _06459_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15229_ clknet_leaf_15_i_clk _00774_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07982_ _01579_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__xnor2_1
X_09721_ _03124_ _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09652_ _03063_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__nor2_1
X_08603_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _02134_
+ _02135_ _02055_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__o221a_1
X_09583_ _02988_ _02996_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08534_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\] _02072_ VGND VGND VPWR
+ VPWR _02073_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08465_ _01879_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07416_ _01095_ net249 _01150_ _01151_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08396_ _01946_ _01948_ _01882_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07347_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _01077_ VGND
+ VGND VPWR VPWR _01090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07278_ _01021_ _01022_ _01023_ _01024_ _01026_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09017_ _02498_ _02493_ _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold150 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold194 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _03295_ VGND
+ VGND VPWR VPWR _03296_ sky130_fd_sc_hd__xnor2_1
X_12930_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05912_
+ _05845_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__o21ai_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _05855_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__nand2_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ clknet_leaf_44_i_clk _00145_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11812_ _04943_ _04947_ _04948_ _04758_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__o31ai_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _05795_ _05796_ _05794_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ clknet_leaf_39_i_clk _00077_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11743_ _04886_ _04887_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__and2_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ clknet_leaf_36_i_clk _00008_ VGND VGND VPWR VPWR r_i_alpha1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11674_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _04825_
+ _04755_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13413_ _06202_ _06330_ _06331_ _06110_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__o211a_1
X_10625_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14393_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _07156_ VGND
+ VGND VPWR VPWR _07175_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10556_ _03855_ _03856_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ _03605_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__a2bb2o_1
X_13344_ _06268_ _06271_ _06201_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10487_ _03787_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__clkbuf_4
X_13275_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15014_ clknet_4_5_0_i_clk _00559_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12226_ _05282_ _05285_ _05296_ _05302_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__or4_4
X_12157_ _05245_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _05246_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_75_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11108_ _04341_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__and2_1
X_12088_ _05153_ net529 _05185_ _05186_ _05170_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__o221a_1
X_11039_ _04272_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14729_ clknet_leaf_73_i_clk _00274_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08250_ _01717_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\] _01823_ _01827_
+ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08181_ net29 net47 VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__xor2_2
XFILLER_0_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07965_ net48 net30 VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__or2b_1
X_09704_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03098_ VGND
+ VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nand2_1
X_07896_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\] _01509_ VGND VGND
+ VPWR VPWR _01510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09635_ _02770_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__nand2_1
X_09566_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02987_ VGND
+ VGND VPWR VPWR _02988_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08517_ _01881_ _02056_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09497_ _02924_ _02913_ _02905_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08448_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\] _01993_ VGND VGND VPWR
+ VPWR _01994_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08379_ _01932_ _01934_ _01882_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10410_ _03703_ _03712_ _03713_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _04375_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04582_
+ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10341_ _03663_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _06003_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__o41ai_2
X_10272_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] _03609_
+ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12011_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04769_ _05125_
+ _05126_ _04965_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13962_ _06292_ net116 VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__nor2_1
X_12913_ _05871_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _05898_ _05899_ _05751_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__o221a_1
X_13893_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND
+ VGND VPWR VPWR _06746_ sky130_fd_sc_hd__or2_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05844_ sky130_fd_sc_hd__clkbuf_4
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05500_ net634 _05495_ _05785_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__o211a_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14514_ clknet_leaf_31_i_clk _00060_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
X_11726_ _04862_ _04871_ _04872_ _04739_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__o211a_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ _07216_ _07219_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__xor2_1
X_11657_ _04769_ net572 _04762_ _04812_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10608_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14376_ _07159_ _07160_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11588_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _04758_
+ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13327_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _06256_ _06257_ _06197_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10539_ _03839_ _03840_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13258_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12209_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05291_ _05282_
+ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__o21ba_1
X_13189_ _06136_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07750_ _01003_ _01395_ net7 VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__o21ai_1
X_07681_ net19 _01347_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09420_ _02844_ net515 _02854_ _02855_ _02827_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09351_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _02797_
+ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08302_ _01867_ net203 _01823_ _01871_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09282_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _02726_ _02733_
+ _02735_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_47_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08233_ _01717_ net309 _01635_ _01813_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08164_ _01750_ _01725_ _01738_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08095_ net42 net24 VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08997_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__or2_1
X_07948_ net39 net21 VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__or2b_1
X_07879_ _01493_ _01494_ _01495_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__a21o_1
X_09618_ _03024_ _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__and2_1
X_10890_ _04135_ _04139_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09549_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR
+ VPWR _02972_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12560_ _05592_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11511_ _04690_ _04061_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_4
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12491_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _05522_
+ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__or2_1
Xwire113 _06051_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_1
X_14230_ _06905_ _07033_ _07034_ _06996_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11442_ _04468_ _04628_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11373_ _04567_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__and2_1
X_14161_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06974_
+ _06904_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13112_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ _05877_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__o21a_1
X_10324_ _03649_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__buf_2
X_14092_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND VPWR
+ VPWR _06917_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _05998_ _06012_ _06013_ _05938_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__o211a_1
X_10255_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03572_ _03596_
+ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__a21o_1
X_10186_ _03207_ _03536_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__nand2_1
X_14994_ clknet_leaf_109_i_clk _00539_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13945_ _06788_ _06789_ _06553_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__o21a_1
X_13876_ _06729_ _06730_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__xnor2_1
X_12827_ _05807_ _05821_ _05817_ _05826_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _04754_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__or2_1
X_12689_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05706_ VGND
+ VGND VPWR VPWR _05707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14428_ _07191_ _07192_ _07200_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14359_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _07144_ VGND
+ VGND VPWR VPWR _07146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08920_ _02152_ net649 _02333_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__a21o_1
X_08851_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02349_
+ _02344_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__o21a_1
X_07802_ net4 net5 _01431_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__and3_2
X_08782_ _02297_ _01549_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _02298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07733_ _01387_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
X_07664_ net202 _01333_ _01336_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_95_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09403_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _02837_
+ _02840_ _02751_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07595_ diff_valid VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09334_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _02776_
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND VPWR
+ VPWR _02783_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09265_ _02117_ _02712_ _01958_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08216_ _01717_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\] _01635_ _01799_
+ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__o211a_1
X_09196_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _02661_ VGND
+ VGND VPWR VPWR _02662_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08147_ _01737_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08078_ _01637_ _01671_ _01651_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10040_ _03389_ _03405_ _03406_ _03292_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__o211a_1
Xhold10 _00429_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _00195_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net105 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 net95 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net101 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold87 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _04850_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__and2_1
Xhold98 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13730_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06599_
+ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__nor2_1
X_10942_ _04179_ _04184_ _04192_ _04188_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13661_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06514_ VGND
+ VGND VPWR VPWR _06549_ sky130_fd_sc_hd__xor2_1
X_10873_ _04096_ _04104_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15400_ clknet_leaf_30_i_clk _00945_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12612_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13592_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06488_ VGND
+ VGND VPWR VPWR _06489_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15331_ clknet_leaf_18_i_clk _00876_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12543_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05577_ VGND
+ VGND VPWR VPWR _05578_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15262_ clknet_leaf_10_i_clk _00807_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12474_ _05500_ net519 _05519_ _05520_ _05391_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14213_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _07018_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__or3b_1
X_11425_ _04611_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__nor2_1
X_15193_ clknet_leaf_0_i_clk _00738_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14144_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _06951_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__and3_1
X_11356_ _04549_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10307_ _03634_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__or2_1
X_14075_ _06903_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__clkbuf_4
X_11287_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04489_ VGND
+ VGND VPWR VPWR _04490_ sky130_fd_sc_hd__xor2_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _05842_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__clkbuf_4
X_10238_ _03574_ _03578_ _03583_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a21bo_1
X_10169_ _03206_ _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_11_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_11_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14977_ clknet_leaf_88_i_clk _00522_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13928_ _06774_ _06775_ _06584_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13859_ _06707_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07380_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _01105_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__or3_4
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09050_ _02524_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08001_ _01599_ _01601_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold502 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold513 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\] VGND VGND VPWR VPWR
+ net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09952_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _03324_ VGND
+ VGND VPWR VPWR _03326_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08903_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _02394_
+ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__or2_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__nand2_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02335_
+ _02337_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__o21ai_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[15\] VGND VGND VPWR VPWR
+ _02282_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_18_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ net11 _01371_ _01344_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__a21o_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08696_ _01866_ _02218_ _02219_ _01552_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07647_ _01323_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07578_ diff1\[3\] diff2\[3\] _01259_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09317_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] _02758_
+ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ _02329_ net534 _02381_ _02709_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09179_ _02322_ net567 _02645_ _02646_ _02414_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11210_ _04420_ _04422_ _04414_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__mux2_1
X_12190_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05260_ VGND
+ VGND VPWR VPWR _05276_ sky130_fd_sc_hd__or2_1
X_11141_ _04364_ _04366_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR out_alpha[17] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 VGND VGND VPWR VPWR out_costheta[10] sky130_fd_sc_hd__clkbuf_4
X_11072_ _04295_ _04303_ _04304_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__a21bo_1
Xoutput88 net88 VGND VGND VPWR VPWR out_costheta[4] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 VGND VGND VPWR VPWR out_sintheta[14] sky130_fd_sc_hd__clkbuf_4
X_14900_ clknet_leaf_87_i_clk _00445_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10023_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__or2_1
X_14831_ clknet_leaf_77_i_clk net604 VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14762_ clknet_leaf_73_i_clk _00307_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_4
X_11974_ _05093_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13713_ _06588_ _06589_ _06590_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__a21oi_1
X_10925_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04177_ VGND
+ VGND VPWR VPWR _04178_ sky130_fd_sc_hd__xnor2_1
X_14693_ clknet_leaf_57_i_clk _00238_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13644_ _06534_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
X_10856_ _04097_ _04114_ _04103_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _06454_ _06464_ _06465_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__o21ai_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04049_
+ _04035_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__o21a_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ clknet_leaf_22_i_clk _00859_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _05488_ _05563_ _05564_ _05343_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15245_ clknet_leaf_10_i_clk _00790_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12457_ _05500_ net552 _05505_ _05506_ _05391_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11408_ _04592_ _04594_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__a21oi_1
X_15176_ clknet_leaf_114_i_clk _00721_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12388_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05423_ VGND
+ VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14127_ _06646_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__nor2_1
X_11339_ _01251_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14058_ _06839_ _06864_ _06885_ _06889_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__and4_1
X_13009_ _05978_ _05979_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__o21ai_1
X_08550_ _02086_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07501_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _01045_ _01013_
+ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__o21a_1
X_08481_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR VPWR
+ _02024_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07432_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _01154_ VGND
+ VGND VPWR VPWR _01166_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07363_ _01095_ net233 _01103_ _01104_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09102_ net273 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] VGND
+ VGND VPWR VPWR _02577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07294_ _01036_ _01041_ _01026_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09033_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _02514_ VGND
+ VGND VPWR VPWR _02515_ sky130_fd_sc_hd__xor2_2
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold310 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 diff2\[16\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold343 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND VGND VPWR
+ VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold398 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09935_ _03182_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] VGND
+ VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nand2_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _03244_
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND VPWR
+ VPWR _03252_ sky130_fd_sc_hd__a21o_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _01959_ _02324_ _02325_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__and3_1
X_09797_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__or2_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _02263_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__nor2_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _02202_ _02203_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__and2_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__clkbuf_4
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _04835_ VGND
+ VGND VPWR VPWR _04839_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10641_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03933_ VGND
+ VGND VPWR VPWR _03934_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13360_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _06283_ _06284_ _06285_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__o221a_1
X_10572_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03870_ VGND
+ VGND VPWR VPWR _03871_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12311_ _05377_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _05382_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13291_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _06224_
+ _06225_ _06216_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15030_ clknet_leaf_98_i_clk _00575_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12242_ _05310_ _05320_ _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__o21a_1
X_12173_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05236_ VGND VGND
+ VPWR VPWR _05260_ sky130_fd_sc_hd__or4_4
X_11124_ _04356_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
X_11055_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04293_ VGND
+ VGND VPWR VPWR _04294_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10006_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _03375_ sky130_fd_sc_hd__inv_2
X_14814_ clknet_leaf_68_i_clk _00359_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14745_ clknet_leaf_56_i_clk _00290_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11957_ _04862_ _05078_ _05079_ _05080_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10908_ _04162_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14676_ clknet_leaf_57_i_clk _00221_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11888_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05016_ VGND
+ VGND VPWR VPWR _05017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13627_ _06516_ _06519_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10839_ _04011_ net333 _04003_ _04099_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13558_ _04455_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12509_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _05539_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13489_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15228_ clknet_leaf_15_i_clk _00773_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15159_ clknet_leaf_122_i_clk _00704_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07981_ _01565_ _01571_ _01564_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__a21o_1
X_09720_ _03110_ _03115_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09651_ _03051_ _03054_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__nor2_1
X_08602_ _02126_ _02129_ _02133_ _01870_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__o31ai_1
X_09582_ _02988_ _02982_ _02996_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08533_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\] _02071_ VGND VGND VPWR
+ VPWR _02072_ sky130_fd_sc_hd__xor2_2
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08464_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[6\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\]
+ _01992_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07415_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08395_ _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07346_ _01016_ net279 _01087_ _01089_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07277_ _01025_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09016_ _02498_ _02493_ _02486_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold140 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _00325_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 net108 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _00254_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _03295_ sky130_fd_sc_hd__o21ba_1
X_09849_ _03190_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__clkbuf_4
X_12860_ _05844_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__clkbuf_4
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _04943_ _04947_ _04948_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__o21a_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _05799_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ clknet_leaf_39_i_clk _00076_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11742_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04885_ VGND
+ VGND VPWR VPWR _04887_ sky130_fd_sc_hd__or2_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14461_ clknet_leaf_36_i_clk _00007_ VGND VGND VPWR VPWR r_i_alpha1\[11\] sky130_fd_sc_hd__dfxtp_1
X_11673_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _04825_
+ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__nor2_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13412_ _06251_ net512 VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__or2_1
X_10624_ _03626_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03917_
+ _03918_ _03814_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14392_ _06910_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _01766_
+ _07174_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13343_ _06269_ _06270_ _06235_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10555_ _03852_ _03854_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13274_ _06210_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ _06203_ _06212_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10486_ _03623_ _03794_ _03795_ _03780_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__o211a_1
X_15013_ clknet_leaf_90_i_clk _00558_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12225_ _05305_ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__nand2_1
X_12156_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05244_ VGND
+ VGND VPWR VPWR _05245_ sky130_fd_sc_hd__xor2_1
X_11107_ _04336_ _04340_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__or2_1
X_12087_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _05184_
+ _01250_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__o21ai_1
X_11038_ _04064_ _04271_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12989_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _05963_ VGND
+ VGND VPWR VPWR _05965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14728_ clknet_leaf_72_i_clk _00273_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14659_ clknet_leaf_54_i_clk _00204_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08180_ _01749_ _01754_ _01768_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07964_ _01565_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09703_ _03090_ _03099_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07895_ _01329_ _01507_ _01503_ _01508_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__a22oi_2
X_09634_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__or4_2
X_09565_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _02984_ _02986_
+ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_78_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08516_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\]
+ _02034_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__or3_1
X_09496_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR _02924_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08447_ _01880_ _01992_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08378_ _01933_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07329_ _01068_ _01073_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10340_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _03657_
+ _03651_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10271_ _03607_ net132 _03568_ _03611_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__o211a_1
X_12010_ _05116_ _05120_ _05124_ _04754_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__a31o_1
X_13961_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__nor4_1
X_12912_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05897_
+ _05845_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__o21ai_1
X_13892_ _06743_ _06744_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__xnor2_1
X_12843_ _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__clkbuf_4
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _05783_ _05784_ _05501_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__o21ai_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ clknet_leaf_31_i_clk _00059_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_1
X_11725_ _04765_ net497 VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__or2_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14444_ _07018_ _07157_ _07195_ _07204_ _07218_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11656_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _04810_
+ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10607_ _03899_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14375_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _07144_ VGND
+ VGND VPWR VPWR _07160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11587_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13326_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06255_
+ _06232_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10538_ _03836_ _03838_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13257_ _06199_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__clkbuf_4
X_10469_ _01474_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12208_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05291_ _05286_
+ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13188_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06136_ VGND
+ VGND VPWR VPWR _06141_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12139_ _05215_ _05219_ _05216_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07680_ net19 _01347_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09350_ _02795_ _02796_ _02772_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08301_ net155 _01870_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09281_ _02739_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08232_ _01330_ _01642_ _01811_ _01812_ _01485_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08163_ net27 net45 _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08094_ _01539_ net632 _01685_ _01688_ _01661_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08996_ _02465_ _02478_ _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__a21o_1
X_07947_ net21 net39 VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07878_ _01493_ _01494_ _01464_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__o21ai_1
X_09617_ _02750_ _03029_ _03030_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__a31o_1
X_09548_ _02748_ _02970_ _02971_ _02260_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09479_ _02907_ _02898_ _02901_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__o31a_1
XFILLER_0_93_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11510_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ _04671_ _04412_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__o31a_1
XFILLER_0_108_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12490_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _05528_
+ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11441_ _04626_ _04627_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ _04375_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_136_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14160_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06974_
+ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__nor2_1
X_11372_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04565_ VGND
+ VGND VPWR VPWR _04568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13111_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _06071_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10323_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _03649_ sky130_fd_sc_hd__inv_2
X_14091_ _06910_ net318 _06915_ _06916_ _06631_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13042_ _05848_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND
+ VGND VPWR VPWR _06013_ sky130_fd_sc_hd__or2_1
X_10254_ _03591_ _03598_ _02132_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10185_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _03521_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__or3_4
X_14993_ clknet_leaf_108_i_clk _00538_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13944_ _06788_ _06789_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__nand2_1
X_13875_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _06716_ _06726_
+ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__a21o_1
X_12826_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05789_ VGND
+ VGND VPWR VPWR _05829_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12757_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__or2_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _04844_ _04846_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_72_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12688_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14427_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _07157_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__o21a_1
X_11639_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _04778_ _04795_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14358_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _07144_ VGND
+ VGND VPWR VPWR _07145_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13309_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _06228_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14289_ _07077_ _07081_ _07076_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08850_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02348_
+ _02344_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07801_ net198 _01345_ _01433_ _01434_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__a22o_1
X_08781_ _01549_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__nor2_1
X_07732_ net379 _01386_ _01358_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07663_ _00991_ _01334_ _01335_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__a21oi_1
X_09402_ _02837_ _02840_ net267 VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07594_ r_i_alpha1\[5\] _01280_ _01276_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__mux2_1
X_09333_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02777_
+ _02409_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09264_ _02710_ _02724_ _02132_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08215_ _01465_ _01798_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09195_ _02520_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__xnor2_1
X_08146_ _01735_ _01736_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__and2b_1
X_08077_ _01638_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND VGND
+ VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 _00599_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 _00709_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _02457_ _02460_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__o21ai_1
Xhold55 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 diff2\[11\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05108_ _04757_
+ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__mux2_1
Xhold88 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13660_ _06548_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
X_10872_ _04113_ _04123_ _04114_ _04103_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12611_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05526_ _05639_
+ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__a21o_1
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13591_ _06463_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15330_ clknet_leaf_18_i_clk _00875_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_12542_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ _05525_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15261_ clknet_leaf_10_i_clk _00806_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12473_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05518_
+ _05490_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14212_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__or2_1
X_11424_ _04233_ _04610_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__nor2_1
X_15192_ clknet_leaf_0_i_clk _00737_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14143_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _06946_ VGND VGND
+ VPWR VPWR _06960_ sky130_fd_sc_hd__or4_1
X_11355_ _04529_ _04535_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10306_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND VPWR
+ VPWR _03635_ sky130_fd_sc_hd__a21oi_1
X_14074_ _06902_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__clkbuf_4
X_11286_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04481_ _04413_
+ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _05843_ _05996_ _05997_ _05938_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__o211a_1
X_10237_ _03583_ _03578_ _03574_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__and3b_1
X_10168_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _03477_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__or4_4
X_14976_ clknet_leaf_90_i_clk _00521_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_10099_ _03456_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13927_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__nor2_1
X_13858_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _06707_ VGND
+ VGND VPWR VPWR _06715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12809_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND
+ VGND VPWR VPWR _05815_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13789_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06653_ VGND
+ VGND VPWR VPWR _06654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08000_ _01589_ _01591_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold503 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR VPWR
+ net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR
+ VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09951_ _03324_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _03325_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08902_ _02321_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _02381_ _02398_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03260_
+ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__nor2_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _02329_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _02338_ _02339_ _02309_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08764_ _02281_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
X_07715_ net11 _01371_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__nor2_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _01873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _02219_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07646_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[15\] _01322_ diff_valid
+ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07577_ _01266_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09316_ _02757_ net313 _02766_ _02767_ _02689_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09247_ _02705_ _02707_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09178_ _02638_ _02631_ _02644_ _02369_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08129_ _01719_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11140_ _04164_ _04338_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput67 net67 VGND VGND VPWR VPWR out_alpha[1] sky130_fd_sc_hd__clkbuf_4
X_11071_ _04012_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04307_
+ _04308_ _04059_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__o221a_1
Xoutput78 net78 VGND VGND VPWR VPWR out_costheta[11] sky130_fd_sc_hd__clkbuf_4
Xoutput89 net89 VGND VGND VPWR VPWR out_costheta[5] sky130_fd_sc_hd__clkbuf_4
X_10022_ _03183_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__clkbuf_4
X_14830_ clknet_leaf_77_i_clk _00375_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11973_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05072_ VGND
+ VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nand2_1
X_14761_ clknet_leaf_72_i_clk _00306_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10924_ _04166_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__clkbuf_4
X_13712_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR _06590_ sky130_fd_sc_hd__inv_2
X_14692_ clknet_leaf_57_i_clk _00237_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10855_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04095_ _04102_
+ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__a21bo_1
X_13643_ _06501_ _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__and2_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13574_ _06456_ _06466_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__or2_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _04048_ _04052_ _04053_ _03780_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__o211a_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _05492_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__or2_1
X_15313_ clknet_leaf_23_i_clk _00858_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12456_ _05203_ _05503_ _05504_ _05487_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__a31o_1
X_15244_ clknet_leaf_11_i_clk _00789_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11407_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _04545_ VGND
+ VGND VPWR VPWR _04598_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15175_ clknet_leaf_114_i_clk _00720_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12387_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05423_ VGND
+ VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14126_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _06941_
+ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__or2_1
X_11338_ _04521_ _04530_ _04535_ _04396_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14057_ _06878_ _06879_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__nor2_1
X_11269_ _04462_ _04464_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__nand2_1
X_13008_ _05979_ _05980_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_118_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14959_ clknet_leaf_90_i_clk _00504_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_07500_ _01076_ _01148_ _01145_ _01080_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__a221o_1
X_08480_ _02014_ _02018_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__nand2_1
X_07431_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _01154_ VGND
+ VGND VPWR VPWR _01165_ sky130_fd_sc_hd__nor2_2
Xclkbuf_4_9_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_9_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07362_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__o21a_1
X_09101_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07293_ _01037_ _01040_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09032_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _02504_ _02343_
+ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold300 net71 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold322 net85 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 diff1\[0\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold344 _00549_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 diff2\[14\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 net79 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net516 sky130_fd_sc_hd__buf_1
X_09934_ _03298_ _03300_ _03308_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09865_ _03249_ _03250_ _02851_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__a21oi_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nand2_1
X_09796_ net141 _03189_ _03017_ _03192_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08747_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\] _02264_ _02265_ VGND
+ VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21o_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\] _02201_ VGND VGND VPWR
+ VPWR _02203_ sky130_fd_sc_hd__or2_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ diff2\[12\] _01270_ _01272_ diff3\[12\] _01308_ VGND VGND VPWR VPWR _01309_
+ sky130_fd_sc_hd__a221o_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03920_ _03650_
+ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10571_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _03862_ _03649_
+ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12310_ _05140_ net289 _05141_ _05381_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13290_ _06224_ _06225_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12241_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _05291_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12172_ _05259_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11123_ _03976_ _04355_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__and2_1
X_11054_ _04192_ net115 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_64_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10005_ _03367_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__inv_2
X_14813_ clknet_leaf_68_i_clk _00358_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_79_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14744_ clknet_leaf_73_i_clk _00289_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11956_ _04455_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10907_ _03976_ _04161_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11887_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05015_
+ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__nor2_1
X_14675_ clknet_leaf_57_i_clk _00220_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10838_ _04097_ _04098_ _04012_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o21ai_1
X_13626_ _06492_ _06517_ _06518_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_144_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10769_ _04036_ _04037_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13557_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _06458_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12508_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05535_ VGND VGND
+ VPWR VPWR _05549_ sky130_fd_sc_hd__or4_1
X_13488_ _06352_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15227_ clknet_leaf_111_i_clk _00772_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_12439_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] _05492_
+ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_17_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15158_ clknet_leaf_122_i_clk _00703_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14109_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _06931_
+ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__and2_1
X_15089_ clknet_leaf_120_i_clk _00634_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_07980_ _01562_ _01582_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09650_ _03061_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__nor2_2
X_08601_ _02126_ _02129_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__o21a_1
X_09581_ _02999_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08532_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\] _02056_ _01880_ VGND
+ VGND VPWR VPWR _02071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08463_ _01891_ net608 _02006_ _02007_ _01908_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07414_ _01076_ _01145_ _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__a21o_1
X_08394_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] _01933_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[14\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND VPWR VPWR _01947_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07345_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07276_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09015_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _02498_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 diff3\[6\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 net92 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _03284_ _03288_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nor2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ net252 _03189_ _03235_ _03236_ _03013_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__o221a_1
X_09779_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _02804_ VGND
+ VGND VPWR VPWR _03180_ sky130_fd_sc_hd__or2_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04930_ VGND
+ VGND VPWR VPWR _04948_ sky130_fd_sc_hd__xnor2_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05652_ _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__and2_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04885_ VGND
+ VGND VPWR VPWR _04886_ sky130_fd_sc_hd__nand2_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _04823_ _04824_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__or2b_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ clknet_leaf_40_i_clk _00006_ VGND VGND VPWR VPWR r_i_alpha1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10623_ _03915_ _03916_ _03631_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13411_ _06323_ _06329_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14391_ _07172_ _07173_ _06911_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13342_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06262_
+ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__nor2_1
X_10554_ _03852_ _03854_ _03605_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13273_ _06211_ net456 VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__nand2_1
X_10485_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _03795_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15012_ clknet_leaf_103_i_clk _00557_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12224_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05279_ VGND
+ VGND VPWR VPWR _05306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12155_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] net121 _05163_
+ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__o21a_1
X_11106_ _04336_ _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__nand2_1
X_12086_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _05184_
+ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__and2_1
X_11037_ _04277_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
X_12988_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _05963_ VGND
+ VGND VPWR VPWR _05964_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14727_ clknet_leaf_73_i_clk _00272_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11939_ _05062_ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14658_ clknet_leaf_45_i_clk _00203_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13609_ _06502_ _06503_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__and2_1
X_14589_ clknet_leaf_37_i_clk _00134_ VGND VGND VPWR VPWR diff3\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07963_ net21 net39 _01557_ _01566_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09702_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _03109_ VGND
+ VGND VPWR VPWR _03110_ sky130_fd_sc_hd__xor2_2
XFILLER_0_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07894_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\] _01502_ VGND VGND
+ VPWR VPWR _01508_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09633_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _03047_ sky130_fd_sc_hd__inv_2
X_09564_ _02985_ _02771_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__mux2_2
XFILLER_0_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08515_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _02053_
+ _02054_ _02055_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09495_ _02921_ _02922_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__and2_1
X_08446_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[4\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[3\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\]
+ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__or4_2
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08377_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[11\] _01928_ VGND VGND
+ VPWR VPWR _01933_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07328_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _01017_ _01052_
+ _01071_ _01072_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07259_ _01009_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10270_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _03609_
+ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13960_ _06798_ _06800_ _06797_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__a21o_1
X_12911_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05897_
+ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__and2_1
X_13891_ _06736_ _06740_ _06734_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__o21ai_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__clkbuf_4
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05782_ _05779_ _05780_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__and3_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ clknet_leaf_31_i_clk _00058_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_1
X_11724_ _04863_ _04870_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__xor2_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11655_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _04810_
+ _04770_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__o21ai_1
X_14443_ _07172_ _07194_ _07217_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10606_ _03860_ _03884_ _03901_ _03893_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__or4_1
X_11586_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _04757_ sky130_fd_sc_hd__clkbuf_4
X_14374_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _07144_ VGND
+ VGND VPWR VPWR _07159_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10537_ _03836_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__and2_1
X_13325_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06255_
+ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10468_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND
+ VGND VPWR VPWR _03779_ sky130_fd_sc_hd__or2_1
X_13256_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _06199_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12207_ _05279_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__clkbuf_4
X_13187_ _05854_ net494 _05847_ _06140_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__o211a_1
X_10399_ _03699_ _03715_ _03703_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12138_ _05227_ _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__and2b_1
X_12069_ _05153_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _05168_ _05169_ _05170_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08300_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09280_ _02738_ _01979_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08231_ _01638_ _01810_ _01472_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08162_ _01741_ _01751_ _01738_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08093_ _01556_ _01687_ _01480_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08995_ _02465_ _02460_ _02475_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__a31o_1
X_07946_ _01454_ _01548_ _01551_ _01552_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07877_ _01488_ _01490_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] VGND
+ VGND VPWR VPWR _01494_ sky130_fd_sc_hd__mux2_1
X_09616_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out _03031_ VGND
+ VGND VPWR VPWR _03032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09547_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _02971_ sky130_fd_sc_hd__or2_1
X_09478_ _02898_ _02901_ _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08429_ _01969_ _01970_ _01975_ _01868_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__o31a_1
XFILLER_0_108_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11440_ _04623_ _04625_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__nor2_1
Xwire115 _04269_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_1
XFILLER_0_135_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11371_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04565_ VGND
+ VGND VPWR VPWR _04567_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13110_ _06064_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _06070_ sky130_fd_sc_hd__and2b_1
X_10322_ _03625_ net501 _03647_ _03648_ _03633_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14090_ _06647_ _06913_ _06914_ _06904_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13041_ _06009_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10253_ _03596_ _03597_ _03186_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10184_ _01765_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14992_ clknet_leaf_108_i_clk _00537_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13943_ _06774_ _06781_ _06780_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13874_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _06707_ VGND
+ VGND VPWR VPWR _06729_ sky130_fd_sc_hd__xnor2_1
X_12825_ _05501_ net563 _05827_ _05828_ _05751_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _05767_ VGND
+ VGND VPWR VPWR _05768_ sky130_fd_sc_hd__and2_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11707_ _04853_ _04854_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__nor2_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _05500_ net315 _05495_ _05705_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14426_ _07059_ net451 VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__nand2_1
X_11638_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _04789_
+ _04795_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14357_ _07135_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__clkbuf_4
X_11569_ _04728_ _04722_ _04731_ _04735_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13308_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _06218_ VGND VGND
+ VPWR VPWR _06241_ sky130_fd_sc_hd__and4_1
X_14288_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _07041_ VGND
+ VGND VPWR VPWR _07084_ sky130_fd_sc_hd__xnor2_1
X_13239_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06142_ VGND
+ VGND VPWR VPWR _06185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07800_ net4 _01431_ _00993_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__o21a_1
X_08780_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[16\] _02283_ VGND VGND VPWR
+ VPWR _02296_ sky130_fd_sc_hd__nor2_2
X_07731_ _01384_ _01385_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07662_ _00991_ _01334_ _00992_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09401_ _02409_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__xor2_1
X_07593_ diff2\[5\] _01270_ _01272_ diff3\[5\] _01279_ VGND VGND VPWR VPWR _01280_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09332_ _02757_ net495 _02780_ _02781_ _02689_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09263_ _02722_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08214_ _01602_ _01797_ _01329_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09194_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02652_ _02342_
+ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08145_ net45 net27 VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08076_ _01670_ _01671_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 _00594_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _02463_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__and2_1
Xhold45 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _00487_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 _00650_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[14\] _01536_
+ _01538_ _01513_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__o221a_1
Xhold78 diff2\[9\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 CORDIC_PE\[0\].genblk1.cordic_engine_inst.i_quadrant\[0\] VGND VGND VPWR VPWR
+ net206 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ _04189_ _04190_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10871_ _04111_ _04121_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12610_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05625_ VGND
+ VGND VPWR VPWR _05639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13590_ _06450_ _06472_ _06473_ _06481_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__or4_2
XFILLER_0_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12541_ _05488_ _05575_ _05576_ _05343_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15260_ clknet_leaf_10_i_clk _00805_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12472_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05518_
+ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14211_ _06904_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] VGND
+ VGND VPWR VPWR _07017_ sky130_fd_sc_hd__and2_1
X_11423_ _04233_ _04610_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__and2_1
X_15191_ clknet_leaf_0_i_clk _00736_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11354_ _04550_ _04534_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__a21oi_1
X_14142_ _06928_ net346 _06958_ _06959_ _06922_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10305_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND VPWR
+ VPWR _03634_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11285_ _04442_ _04487_ _04488_ _04456_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__o211a_1
X_14073_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _06902_ sky130_fd_sc_hd__inv_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13024_ _05848_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _05997_ sky130_fd_sc_hd__or2_1
X_10236_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03572_ VGND
+ VGND VPWR VPWR _03583_ sky130_fd_sc_hd__xnor2_1
X_10167_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__or2_1
X_14975_ clknet_leaf_93_i_clk _00520_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10098_ _03031_ _03455_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13926_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13857_ _06556_ _06713_ _06714_ _06459_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__o211a_1
X_12808_ _05812_ _05813_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13788_ _06292_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND
+ VGND VPWR VPWR _06653_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _05739_ _05748_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14409_ _07182_ _07184_ _07188_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15389_ clknet_leaf_19_i_clk _00934_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold504 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND VGND VPWR
+ VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold515 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR VPWR
+ net632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold526 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09950_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03323_ VGND
+ VGND VPWR VPWR _03324_ sky130_fd_sc_hd__xor2_1
Xclkbuf_4_5_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_5_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_08901_ _02392_ _02396_ _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__o21ai_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR _03264_ sky130_fd_sc_hd__inv_2
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02336_
+ _02337_ _02333_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__a31o_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _01981_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__and2_1
X_07714_ _01374_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08694_ _02213_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07645_ r_i_alpha1\[15\] _01321_ _01258_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07576_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\] net380 _01255_ VGND
+ VGND VPWR VPWR _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09315_ _02760_ _02765_ _02747_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09246_ _02705_ _02707_ _02319_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09177_ _02638_ _02631_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08128_ _01718_ net44 VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08059_ _01653_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11070_ _04305_ _04306_ _03994_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__a21o_1
Xoutput57 net57 VGND VGND VPWR VPWR o_valid_out sky130_fd_sc_hd__clkbuf_4
Xoutput68 net68 VGND VGND VPWR VPWR out_alpha[2] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 VGND VGND VPWR VPWR out_costheta[12] sky130_fd_sc_hd__clkbuf_4
X_10021_ _03191_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03387_
+ _03388_ _03258_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o221a_1
X_14760_ clknet_leaf_72_i_clk _00305_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_11972_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05072_ VGND
+ VGND VPWR VPWR _05093_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13711_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _06571_ _06587_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__a31o_1
X_10923_ _04153_ _04168_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__or2b_1
X_14691_ clknet_leaf_57_i_clk _00236_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13642_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06532_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__mux2_1
X_10854_ _04111_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _06470_ _06471_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10785_ _03999_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15312_ clknet_leaf_23_i_clk _00857_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05562_
+ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15243_ clknet_leaf_12_i_clk _00788_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12455_ _05503_ _05504_ _05203_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11406_ _04597_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__clkbuf_1
X_15174_ clknet_leaf_114_i_clk _00719_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12386_ _05434_ _05448_ _05449_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14125_ _06910_ net215 _06678_ _06945_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__o211a_1
X_11337_ _04521_ _04530_ _04535_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14056_ _06569_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] VGND
+ VGND VPWR VPWR _06888_ sky130_fd_sc_hd__and2_1
X_11268_ _04471_ _04472_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ _05978_ _05878_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__nor2_1
X_10219_ _03389_ _03566_ _03567_ _03515_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11199_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__buf_2
X_14958_ clknet_leaf_90_i_clk _00503_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13909_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06716_ VGND
+ VGND VPWR VPWR _06759_ sky130_fd_sc_hd__or2_1
X_14889_ clknet_leaf_109_i_clk _00434_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_07430_ _01019_ _01163_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07361_ _01098_ _01102_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09100_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _02574_
+ _02575_ _02414_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07292_ _01038_ _01039_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09031_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02506_ VGND
+ VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold301 diff2\[13\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND VPWR
+ VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold323 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net440 sky130_fd_sc_hd__buf_1
Xhold334 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND VGND
+ VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold345 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _03298_ _03300_ _03308_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _03243_
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND VPWR
+ VPWR _03250_ sky130_fd_sc_hd__o21ai_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__or2_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _03191_ net305 VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08746_ _02252_ _02257_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__and2b_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\] _02201_ VGND VGND VPWR
+ VPWR _02202_ sky130_fd_sc_hd__nand2_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _01273_ diff1\[12\] VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07559_ _01254_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10570_ _03623_ _03868_ _03869_ _03780_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09229_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02685_ _02674_
+ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_90_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12240_ _05307_ _05313_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _04850_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11122_ _04047_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04353_
+ _04354_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__a22o_1
X_11053_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR _04292_ sky130_fd_sc_hd__inv_2
X_10004_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03372_ VGND
+ VGND VPWR VPWR _03373_ sky130_fd_sc_hd__xor2_1
Xclkbuf_0_i_clk i_clk VGND VGND VPWR VPWR clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_14812_ clknet_leaf_67_i_clk _00357_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14743_ clknet_leaf_65_i_clk _00288_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11955_ _04770_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _05079_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10906_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04160_ _03996_
+ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__mux2_1
X_14674_ clknet_leaf_57_i_clk _00219_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_11886_ _04557_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND VGND VPWR VPWR
+ _05015_ sky130_fd_sc_hd__nor4_1
XFILLER_0_39_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13625_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _06514_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__o41ai_2
XFILLER_0_7_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10837_ _04085_ _04092_ _04096_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13556_ _06450_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__xor2_1
X_10768_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR _04038_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12507_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05547_ _05548_ _05544_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13487_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06351_ VGND
+ VGND VPWR VPWR _06396_ sky130_fd_sc_hd__xnor2_1
X_10699_ _03976_ _03986_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15226_ clknet_leaf_111_i_clk _00771_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_12438_ _05488_ net244 _05141_ _05493_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15157_ clknet_leaf_122_i_clk _00702_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_140_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12369_ _05139_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _05436_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14108_ _06929_ _06930_ _06646_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__mux2_1
X_15088_ clknet_leaf_120_i_clk _00633_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14039_ _06862_ _06869_ _06872_ _06569_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08600_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[17\] _02124_ VGND VGND VPWR
+ VPWR _02133_ sky130_fd_sc_hd__xor2_1
X_09580_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _02986_ VGND
+ VGND VPWR VPWR _03000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08531_ _02070_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08462_ _01995_ _02001_ _02005_ _01924_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07413_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _01051_ _01081_
+ _01148_ _01085_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08393_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] _01932_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[14\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND VPWR VPWR _01946_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07344_ _01012_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07275_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_859 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09014_ _01765_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold120 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold131 diff3\[9\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _00489_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold164 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[1\] VGND VGND VPWR VPWR
+ net292 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold186 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net303 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold197 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _03287_ VGND
+ VGND VPWR VPWR _03293_ sky130_fd_sc_hd__and2_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _03234_
+ _03183_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__a21o_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _03177_ _03178_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__xnor2_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\]
+ _02231_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__or3_2
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04884_ VGND
+ VGND VPWR VPWR _04885_ sky130_fd_sc_hd__xnor2_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04817_
+ _04795_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a21o_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13410_ _06327_ _06328_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10622_ _03915_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nor2_1
X_14390_ _07171_ _07169_ _07170_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__nor3_1
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13341_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06263_
+ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10553_ _03853_ _03843_ _03840_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13272_ _06204_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10484_ _03792_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15011_ clknet_leaf_95_i_clk _00556_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12223_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05279_ VGND
+ VGND VPWR VPWR _05305_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12154_ _05234_ _05242_ _05243_ _05080_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__o211a_1
X_11105_ _04337_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__and2_1
X_12085_ _04829_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _05177_ _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__o31a_1
X_11036_ _03976_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12987_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05962_ VGND
+ VGND VPWR VPWR _05963_ sky130_fd_sc_hd__xor2_1
X_14726_ clknet_leaf_56_i_clk _00271_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11938_ _04831_ _05061_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14657_ clknet_leaf_49_i_clk _00202_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11869_ _04999_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13608_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06488_ VGND
+ VGND VPWR VPWR _06503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14588_ clknet_leaf_34_i_clk _00133_ VGND VGND VPWR VPWR diff3\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13539_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06235_ VGND VGND
+ VPWR VPWR _06441_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15209_ clknet_leaf_2_i_clk _00754_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07962_ net30 net48 VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09701_ _02972_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07893_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\] VGND VGND VPWR VPWR
+ _01507_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09632_ _03046_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09563_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _02984_
+ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__or2_1
X_08514_ _01512_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09494_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02920_ VGND
+ VGND VPWR VPWR _02922_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08445_ _01974_ _01976_ _01986_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08376_ _01926_ _01927_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07327_ _01056_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07258_ net178 net11 _01000_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12910_ _05567_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _05890_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__o31a_1
X_13890_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06707_ VGND
+ VGND VPWR VPWR _06743_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12841_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05841_ sky130_fd_sc_hd__inv_2
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ _05779_ _05780_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__a21oi_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ clknet_leaf_31_i_clk _00057_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11723_ _04868_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__nor2_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _07209_ _07205_ _07213_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__and3_1
X_11654_ _04445_ _04807_ _04809_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10605_ _03867_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14373_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ _07157_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11585_ _04755_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13324_ _05928_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _06247_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__o31a_1
XFILLER_0_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10536_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _03837_ VGND
+ VGND VPWR VPWR _03838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13255_ _06198_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10467_ _03776_ _03777_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12206_ _01252_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__buf_2
X_13186_ _06138_ _06139_ _05855_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__o21ai_1
X_10398_ _03705_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__inv_2
X_12137_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05226_ VGND
+ VGND VPWR VPWR _05228_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12068_ _04538_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__clkbuf_4
X_11019_ _04011_ net571 _04219_ _04261_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14709_ clknet_leaf_51_i_clk net301 VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08230_ _01638_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08161_ _01722_ _01724_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08092_ _01681_ _01686_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08994_ _02463_ _02472_ _02474_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07945_ _01455_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__buf_4
X_07876_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[7\] VGND VGND VPWR VPWR
+ _01493_ sky130_fd_sc_hd__inv_2
X_09615_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _03031_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09546_ _02962_ _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__xnor2_1
X_09477_ _02905_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08428_ _01969_ _01970_ _01975_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire116 _06805_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08359_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND VPWR VPWR
+ _01918_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11370_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04565_ _04552_
+ _04562_ _04547_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10321_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03646_
+ _03642_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__o21ai_1
X_13040_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _06010_ _06005_
+ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__a21o_1
X_10252_ _03595_ _03593_ _03594_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__or3_1
X_10183_ _03191_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03533_
+ _03534_ _03258_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__o221a_1
X_14991_ clknet_leaf_109_i_clk _00536_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13942_ _06786_ _06787_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__nor2_1
X_13873_ _06728_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
X_12824_ _05820_ _05822_ _05826_ _05486_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12755_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05756_ VGND
+ VGND VPWR VPWR _05767_ sky130_fd_sc_hd__nor2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04852_ VGND
+ VGND VPWR VPWR _04854_ sky130_fd_sc_hd__nor2_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12686_ _05703_ _05704_ _05501_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__o21ai_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14425_ _06911_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _07201_
+ _07202_ _01456_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11637_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14356_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _07136_ VGND
+ VGND VPWR VPWR _07143_ sky130_fd_sc_hd__and2_1
X_11568_ _04740_ _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13307_ _06223_ net595 _06239_ _06240_ _06197_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10519_ _03824_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14287_ _07059_ _07082_ _07083_ _06996_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__o211a_1
X_11499_ _04676_ _04680_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13238_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06142_ VGND
+ VGND VPWR VPWR _06184_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13169_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _06112_ VGND
+ VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nand2_1
X_07730_ net18 _01341_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07661_ net14 VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_4
X_09400_ _02757_ net601 _02838_ _02839_ _02827_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07592_ _01273_ diff1\[5\] VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_1_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_09331_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02779_
+ _02755_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09262_ _02717_ _02721_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08213_ _01599_ _01796_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09193_ _02314_ _02658_ _02659_ _02260_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08144_ net27 net45 VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08075_ net38 net56 VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold13 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02462_ VGND
+ VGND VPWR VPWR _02464_ sky130_fd_sc_hd__or2_1
Xhold35 _00596_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _00654_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _01532_ _01537_ _01485_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__o21ai_1
Xhold68 net109 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 diff2\[5\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07859_ _01471_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__nor2_1
X_10870_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _04120_ VGND
+ VGND VPWR VPWR _04127_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09529_ _02950_ _02946_ _02953_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__a21oi_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12540_ _05492_ net607 VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12471_ _05516_ _05517_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14210_ _07016_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11422_ net120 _04609_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__xnor2_1
X_15190_ clknet_leaf_0_i_clk _00735_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14141_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _06957_
+ _06904_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__a21o_1
X_11353_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04520_ _04534_
+ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10304_ _03625_ net592 _03630_ _03632_ _03633_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__o221a_1
X_14072_ _06901_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11284_ _04444_ net491 VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13023_ _05994_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__xnor2_1
X_10235_ _03201_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND
+ VGND VPWR VPWR _03582_ sky130_fd_sc_hd__and2_1
X_10166_ _03517_ _03518_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__and2_1
X_14974_ clknet_leaf_90_i_clk _00519_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10097_ _03031_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__and2_1
X_13925_ _06555_ _06772_ _06773_ _06747_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13856_ _06557_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _06714_ sky130_fd_sc_hd__or2_1
X_12807_ _05806_ _05809_ _05805_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13787_ _06563_ net600 _06651_ _06652_ _06631_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__o221a_1
X_10999_ _04239_ _04241_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12738_ _05501_ net311 _05749_ _05750_ _05751_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__o221a_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12669_ _05632_ _05689_ _05690_ _05675_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14408_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _07156_ VGND
+ VGND VPWR VPWR _07188_ sky130_fd_sc_hd__xor2_1
X_15388_ clknet_leaf_47_i_clk _00933_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14339_ _07124_ _07126_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold505 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND VGND VPWR
+ VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR
+ VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08900_ _02392_ _02396_ _02333_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09880_ _03237_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _03262_ _03263_ _03258_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__o221a_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _02336_ _02337_ net588 VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _01865_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _02278_
+ _02279_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07713_ net392 _01373_ _01358_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__mux2_1
X_08693_ _02194_ _02214_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07644_ diff2\[15\] _01269_ _01271_ diff3\[15\] _01320_ VGND VGND VPWR VPWR _01321_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07575_ _01265_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09314_ _02760_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09245_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _02706_ _02700_
+ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09176_ _02642_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08127_ _01718_ net44 VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08058_ _01638_ _01641_ _01654_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput58 net58 VGND VGND VPWR VPWR out_alpha[0] sky130_fd_sc_hd__clkbuf_4
Xoutput69 net69 VGND VGND VPWR VPWR out_alpha[3] sky130_fd_sc_hd__clkbuf_4
X_10020_ _03383_ _03379_ _03386_ _03201_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__a31o_1
X_11971_ _05082_ _05083_ _05087_ _05091_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__a31o_1
X_13710_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _06580_
+ _06587_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__o21ai_1
X_10922_ _04158_ _04173_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__or2_1
X_14690_ clknet_leaf_56_i_clk _00235_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13641_ _06529_ _06531_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__xor2_1
X_10853_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04110_ VGND
+ VGND VPWR VPWR _04112_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06463_ VGND
+ VGND VPWR VPWR _06471_ sky130_fd_sc_hd__nand2_1
X_10784_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04051_
+ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__xor2_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ clknet_leaf_23_i_clk _00856_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _05560_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__or2b_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15242_ clknet_leaf_11_i_clk _00787_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12454_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11405_ _04468_ _04596_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__and2_1
X_15173_ clknet_leaf_114_i_clk _00718_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12385_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05423_ VGND VGND VPWR
+ VPWR _05449_ sky130_fd_sc_hd__a31o_1
X_14124_ _06911_ _06944_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__nand2_1
X_11336_ net119 _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__xnor2_2
X_14055_ _06563_ net605 _06886_ _06887_ _06631_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__o221a_1
X_11267_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04470_ VGND
+ VGND VPWR VPWR _04472_ sky130_fd_sc_hd__or2_1
X_13006_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05566_ VGND
+ VGND VPWR VPWR _05980_ sky130_fd_sc_hd__nor2_1
X_10218_ _03190_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _03567_ sky130_fd_sc_hd__or2_1
X_11198_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _04412_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10149_ _03499_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14957_ clknet_leaf_90_i_clk _00502_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13908_ _06555_ _06757_ _06758_ _06747_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14888_ clknet_leaf_109_i_clk net378 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13839_ _06688_ _06697_ _06698_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07360_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _01017_ _01052_
+ _01101_ _01072_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07291_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR VPWR
+ _01039_ sky130_fd_sc_hd__o21ai_1
X_09030_ _02512_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold302 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold313 net64 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold335 net90 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR net463 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold357 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _03306_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold379 _03214_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _03243_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__or3_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _02321_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ _01945_ _02323_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__o211a_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _03190_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08745_ _02251_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__inv_2
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08676_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[8\] _02200_ VGND VGND VPWR
+ VPWR _02201_ sky130_fd_sc_hd__xor2_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _01307_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07558_ _01250_ _01253_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07489_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _01159_ _01208_
+ _01209_ _01030_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09228_ _02655_ _02662_ _02663_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09159_ _02608_ _02627_ _02342_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12170_ _05222_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05256_
+ _05257_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11121_ _04350_ _04352_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11052_ _04280_ _04286_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__o21a_1
X_10003_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03371_ VGND
+ VGND VPWR VPWR _03372_ sky130_fd_sc_hd__xnor2_1
X_14811_ clknet_leaf_67_i_clk _00356_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11954_ _05076_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__xnor2_1
X_14742_ clknet_leaf_65_i_clk _00287_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10905_ _04155_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14673_ clknet_leaf_55_i_clk _00218_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_11885_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _05014_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13624_ _06498_ _06504_ _06510_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__and3_1
X_10836_ _04085_ _04092_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13555_ _06454_ _06455_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__or2_1
X_10767_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _04018_ _04035_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12506_ net615 _05546_ _05487_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13486_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06394_
+ _06395_ _06285_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__o221a_1
X_10698_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03985_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15225_ clknet_leaf_111_i_clk _00770_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12437_ net207 _05492_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15156_ clknet_leaf_123_i_clk _00701_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12368_ _05433_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__xnor2_1
X_14107_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _06917_
+ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11319_ _04413_ _04518_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15087_ clknet_leaf_120_i_clk _00632_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12299_ _05128_ _05369_ _05370_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__o31a_1
X_14038_ _06862_ _06869_ _06872_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08530_ _01981_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__and2_1
X_08461_ _01995_ _02001_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07412_ _01146_ _01147_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08392_ _01455_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_4
X_07343_ _01076_ _01079_ _01086_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07274_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _01010_
+ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _02495_
+ _02496_ _02414_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold110 diff1\[9\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _00707_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 net99 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _01233_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _03184_ _03289_ _03291_ _03292_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__o211a_1
X_09846_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _03234_
+ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__nor2_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _03151_ VGND
+ VGND VPWR VPWR _03178_ sky130_fd_sc_hd__xnor2_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02247_
+ _02248_ _02055_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__o221a_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _02173_ _02177_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__nor2_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04819_
+ _04795_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10621_ _03903_ _03910_ _03908_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13340_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR _06268_ sky130_fd_sc_hd__inv_2
X_10552_ _03836_ _03838_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13271_ _06204_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10483_ _03791_ _03782_ _03784_ _03785_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15010_ clknet_leaf_103_i_clk _00555_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_12222_ _05153_ net570 _05303_ _05304_ _05170_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12153_ _05132_ net482 VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11104_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04338_ VGND
+ VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nand2_1
X_12084_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05182_
+ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__nand2_1
X_11035_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _04275_ _03996_
+ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__mux2_1
X_12986_ _05877_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand2_1
X_14725_ clknet_leaf_53_i_clk _00270_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_11937_ _04831_ _05061_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__nor2_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11868_ _04850_ _04998_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14656_ clknet_leaf_49_i_clk _00201_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10819_ _04081_ _03118_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__and2b_1
X_13607_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06488_ VGND
+ VGND VPWR VPWR _06502_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11799_ _04917_ _04918_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14587_ clknet_leaf_34_i_clk _00132_ VGND VGND VPWR VPWR diff3\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13538_ _06432_ _06440_ _04961_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13469_ _06379_ _06380_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ clknet_leaf_2_i_clk _00753_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15139_ clknet_leaf_125_i_clk _00684_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07961_ _01563_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__nor2_2
X_09700_ _02771_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07892_ _01463_ net500 _01460_ _01506_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _03045_ _01979_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09562_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ _02964_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__nor3_2
X_08513_ _02037_ _02044_ _02052_ _01924_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__a31o_1
X_09493_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02920_ VGND
+ VGND VPWR VPWR _02921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08444_ _01990_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08375_ _01891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _01930_ _01931_ _01908_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__o221a_1
X_07326_ _01069_ _01070_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07257_ _01008_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09829_ _03184_ _03219_ _03220_ _03058_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__o211a_1
X_12840_ _05840_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _05781_ VGND
+ VGND VPWR VPWR _05782_ sky130_fd_sc_hd__xnor2_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04867_ VGND
+ VGND VPWR VPWR _04869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ clknet_leaf_31_i_clk _00056_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11653_ _04445_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__nand2_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _07157_ VGND
+ VGND VPWR VPWR _07216_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _03872_ _03873_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14372_ _07156_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__clkbuf_4
X_11584_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13323_ _05927_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10535_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ _03649_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13254_ _05845_ _01979_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10466_ _03765_ _03769_ _03763_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12205_ _05234_ _05288_ _05289_ _05080_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13185_ _06137_ _06133_ _06135_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__and3_1
X_10397_ _03712_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__or2b_1
X_12136_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05226_ VGND
+ VGND VPWR VPWR _05227_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12067_ _05167_ _05165_ _05166_ _05129_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__a31o_1
X_11018_ _04259_ _04260_ _04048_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12969_ _05939_ _05940_ _05945_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14708_ clknet_leaf_51_i_clk _00253_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14639_ clknet_leaf_60_i_clk _00184_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08160_ _01719_ _01720_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08091_ _01669_ _01675_ _01663_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_141_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08993_ _02433_ _02440_ _02447_ _02453_ _02475_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07944_ _01464_ _01550_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__or2_1
X_07875_ _01467_ net528 _01491_ _01492_ _01475_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__o221a_1
X_09614_ _03025_ _03022_ _03028_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__or3b_1
X_09545_ _02967_ _02968_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09476_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02904_ VGND
+ VGND VPWR VPWR _02906_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08427_ _01973_ _01974_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08358_ _01550_ _01916_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07309_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _01010_
+ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08289_ _01454_ _01856_ _01859_ _01860_ _01766_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__o311a_1
XFILLER_0_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10320_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03646_
+ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10251_ _03593_ _03594_ _03595_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__o21a_1
X_10182_ _03531_ _03532_ _03183_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__a21o_1
X_14990_ clknet_leaf_104_i_clk _00535_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_4
X_13941_ _06431_ _06785_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__nor2_1
X_13872_ _06501_ _06727_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12823_ _05820_ _05822_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12754_ _05766_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11705_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04852_ VGND
+ VGND VPWR VPWR _04853_ sky130_fd_sc_hd__and2_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12685_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__nor2_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11636_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _04794_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14424_ _07192_ _07199_ _07200_ _06926_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11567_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04723_ VGND
+ VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nand2_1
X_14355_ _07142_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10518_ _03535_ _03823_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__and2_1
X_13306_ _06238_ _06236_ _06237_ _06216_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__a31o_1
X_14286_ _06907_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _07083_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11498_ _04678_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13237_ _05855_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06182_
+ _06183_ _05910_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__o221a_1
X_10449_ _03280_ _03760_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13168_ _06103_ _06118_ _06117_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__o21a_1
X_12119_ _05132_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _05212_ sky130_fd_sc_hd__or2_1
X_13099_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07660_ _00993_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07591_ _01278_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09330_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02779_
+ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09261_ _02717_ _02721_ _02313_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08212_ _01589_ _01790_ _01587_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09192_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _02659_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08143_ _01717_ net410 _01635_ _01734_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08074_ net56 net38 VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold14 _00426_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02462_ VGND
+ VGND VPWR VPWR _02463_ sky130_fd_sc_hd__nand2_1
Xhold25 _00424_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND VPWR VPWR
+ net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\] _01535_ VGND VGND
+ VPWR VPWR _01537_ sky130_fd_sc_hd__nand2_1
Xhold69 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ _01476_ _01477_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__or2_1
X_07789_ net425 _01425_ _01411_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09528_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _02952_ VGND
+ VGND VPWR VPWR _02953_ sky130_fd_sc_hd__xnor2_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09459_ _02754_ net527 _02749_ _02890_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12470_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05507_
+ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11421_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ _04412_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14140_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _06957_
+ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__nor2_1
X_11352_ net119 VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10303_ _02308_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__clkbuf_4
X_14071_ _06557_ _01979_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__and2_1
X_11283_ _04480_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__xor2_1
X_13022_ _05986_ _05987_ _05984_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10234_ _03189_ net437 _03568_ _03581_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10165_ _03476_ _03499_ _03500_ _03511_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__or4_1
X_14973_ clknet_leaf_90_i_clk _00518_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10096_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03454_ VGND
+ VGND VPWR VPWR _03455_ sky130_fd_sc_hd__xnor2_1
X_13924_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _06773_ sky130_fd_sc_hd__or2_1
X_13855_ _06708_ _06712_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05781_ VGND
+ VGND VPWR VPWR _05812_ sky130_fd_sc_hd__xor2_1
X_10998_ _04239_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__nor2_1
X_13786_ _06650_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _06569_
+ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _04538_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__buf_4
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12668_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND
+ VGND VPWR VPWR _05690_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14407_ _07187_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
X_11619_ _04778_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__or2_1
X_15387_ clknet_leaf_20_i_clk _00932_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_12599_ _05627_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14338_ _07124_ _07126_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold506 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ _07065_ _07066_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__a21oi_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _01958_ _02330_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _02277_ _02270_ _02272_ _01865_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__a31oi_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _01371_ _01372_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__nand2_1
X_08692_ _02194_ _02190_ _02204_ _02215_ _02203_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__a32o_1
X_07643_ diff2\[17\] diff1\[15\] VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07574_ net292 net360 _01255_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09313_ _02763_ _02764_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09244_ _02697_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09175_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _02640_ VGND
+ VGND VPWR VPWR _02643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08126_ net26 VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08057_ net37 net55 VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__and2_1
Xoutput59 net59 VGND VGND VPWR VPWR out_alpha[10] sky130_fd_sc_hd__clkbuf_4
X_08959_ _02433_ _02440_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__o21a_1
X_11970_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ _05081_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__o21a_1
X_10921_ _04139_ _04145_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__or3_1
X_10852_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04110_ VGND
+ VGND VPWR VPWR _04111_ sky130_fd_sc_hd__nand2_1
X_13640_ _06516_ _06519_ _06523_ _06530_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__a31o_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10783_ _03669_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _04041_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__a31o_1
X_13571_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06463_ VGND
+ VGND VPWR VPWR _06470_ sky130_fd_sc_hd__or2_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15310_ clknet_leaf_23_i_clk _00855_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_12522_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _05550_ _05526_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_836 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15241_ clknet_leaf_114_i_clk _00786_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12453_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11404_ _04375_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04594_
+ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__a22o_1
X_12384_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05423_ VGND VGND VPWR
+ VPWR _05448_ sky130_fd_sc_hd__o31a_1
X_15172_ clknet_leaf_113_i_clk _00717_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11335_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04533_ VGND
+ VGND VPWR VPWR _04534_ sky130_fd_sc_hd__xor2_2
XFILLER_0_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14123_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _06943_
+ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11266_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04470_ VGND
+ VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nand2_1
X_14054_ _06877_ _06884_ _06885_ _06569_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__a31o_1
X_13005_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ _05961_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__or3_2
X_10217_ _03564_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__and2_1
X_11197_ _04390_ net460 _04410_ _04411_ _04360_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__o221a_1
X_10148_ _03476_ _03500_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__o21ai_1
X_14956_ clknet_leaf_90_i_clk _00501_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10079_ _03441_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__clkbuf_1
X_13907_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND
+ VGND VPWR VPWR _06758_ sky130_fd_sc_hd__or2_1
X_14887_ clknet_leaf_109_i_clk _00432_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13838_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _06684_ _06685_
+ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__a21o_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13769_ _06293_ _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07290_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR VPWR
+ _01038_ sky130_fd_sc_hd__or3_4
XFILLER_0_116_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15439_ clknet_leaf_31_i_clk _00984_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold303 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net442 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold336 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _00550_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold358 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR VPWR
+ net475 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _03305_ VGND
+ VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nor2_1
Xhold369 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _03237_ net487 _03247_ _03248_ _03013_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__o221a_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _02322_ net300 VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__nand2_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _03185_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\] _02262_ VGND VGND VPWR
+ VPWR _02263_ sky130_fd_sc_hd__xnor2_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[7\] _02191_ _01879_ VGND
+ VGND VPWR VPWR _02200_ sky130_fd_sc_hd__o21a_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[11\] _01306_ _01282_
+ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07557_ _01252_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07488_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _01122_ _01125_
+ _01047_ _01072_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09227_ _02676_ _02686_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09158_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__or2_1
X_08109_ _01675_ _01700_ _01702_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09089_ _02552_ _02557_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__nand2_1
X_11120_ _04350_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11051_ _04278_ _04284_ _04285_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10002_ _03206_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14810_ clknet_leaf_67_i_clk _00355_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_14741_ clknet_leaf_64_i_clk _00286_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_11953_ _05062_ _05065_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__nor2_1
X_10904_ _04139_ _04145_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__o21ai_1
X_14672_ clknet_leaf_55_i_clk _00217_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_11884_ _05005_ _05009_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13623_ _06513_ _06515_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__and2_1
X_10835_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04095_ VGND
+ VGND VPWR VPWR _04096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13554_ _06451_ _06453_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10766_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _04028_
+ _04035_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12505_ net529 _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10697_ _03979_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__xor2_1
X_13485_ _06392_ _06393_ _06216_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__a21o_1
X_15224_ clknet_leaf_15_i_clk net436 VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12436_ _05489_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15155_ clknet_leaf_123_i_clk _00700_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12367_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _05424_ _05426_
+ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14106_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ _06914_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__or3_1
X_11318_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ _04481_ _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__or4_4
X_15086_ clknet_leaf_118_i_clk _00631_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12298_ _05128_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND
+ VGND VPWR VPWR _05371_ sky130_fd_sc_hd__nand2_1
X_11249_ _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__clkbuf_4
X_14037_ _06870_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14939_ clknet_leaf_110_i_clk _00484_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08460_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\] _02004_ VGND VGND VPWR
+ VPWR _02005_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07411_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _01132_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08391_ _01876_ net481 _01823_ _01944_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07342_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _01080_ _01081_
+ _01084_ _01085_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07273_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09012_ _02486_ _02490_ _02494_ _02369_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold100 _00422_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold111 diff1\[5\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 diff2\[10\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[0\] VGND VGND VPWR VPWR
+ net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold177 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _01474_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__clkbuf_4
Xhold199 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _03232_ _03233_ _02850_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__mux2_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03151_ _03174_
+ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__a21o_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _02241_ _02235_ _02246_ _01865_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__a31o_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _02183_ _02184_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__and2b_1
XFILLER_0_139_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ diff2\[8\] _01270_ _01272_ diff3\[8\] _01292_ VGND VGND VPWR VPWR _01293_
+ sky130_fd_sc_hd__a221o_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _01549_ _02122_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nor2_1
X_10620_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03914_ VGND
+ VGND VPWR VPWR _03915_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10551_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10482_ _03782_ _03784_ _03785_ _03791_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__a31oi_4
X_13270_ _06202_ net287 _06203_ _06209_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12221_ _05295_ _05299_ _05302_ _01250_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12152_ _05235_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11103_ _04325_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__clkbuf_4
X_12083_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _05171_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11034_ _04272_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12985_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__or4_1
XFILLER_0_86_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14724_ clknet_leaf_55_i_clk _00269_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11936_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05060_ VGND
+ VGND VPWR VPWR _05061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14655_ clknet_leaf_49_i_clk _00200_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _04770_ _04994_ _04995_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__a31o_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ _01252_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10818_ _04047_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04079_
+ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14586_ clknet_leaf_34_i_clk _00131_ VGND VGND VPWR VPWR diff3\[11\] sky130_fd_sc_hd__dfxtp_1
X_11798_ _04907_ _04918_ _04925_ _04936_ _04926_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_28_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13537_ _06437_ _06438_ _06439_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__a21oi_1
X_10749_ _04016_ _04020_ _03994_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13468_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _06352_ _06376_
+ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15207_ clknet_leaf_1_i_clk _00752_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12419_ _05222_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05477_
+ _05478_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__a22o_1
X_13399_ _06305_ _06309_ _06306_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15138_ clknet_leaf_125_i_clk _00683_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15069_ clknet_leaf_117_i_clk _00614_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_07960_ net31 net49 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__and2b_1
X_07891_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\] _01504_ _01505_ VGND
+ VGND VPWR VPWR _01506_ sky130_fd_sc_hd__a21o_1
X_09630_ _02750_ _03035_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09561_ _02962_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08512_ _02037_ _02044_ _02052_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__a21oi_1
X_09492_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02919_ VGND
+ VGND VPWR VPWR _02920_ sky130_fd_sc_hd__xor2_1
X_08443_ _01981_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08374_ _01926_ _01929_ _01877_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07325_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _01053_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07256_ net376 net10 _01000_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09828_ net126 _03190_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__or2_1
X_09759_ _03152_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND
+ VGND VPWR VPWR _03162_ sky130_fd_sc_hd__and2b_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _05771_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__clkbuf_4
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04867_ VGND
+ VGND VPWR VPWR _04868_ sky130_fd_sc_hd__and2_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _06911_ net518 _07214_ _07215_ _01456_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__o221a_1
X_11652_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _04801_
+ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__and2_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10603_ _03884_ _03897_ _03893_ _03898_ _03892_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__o32a_1
XFILLER_0_92_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14371_ _07144_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11583_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _04754_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13322_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _06241_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10534_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _03836_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13253_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05854_ _06195_
+ _06196_ _06197_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__o221a_1
X_10465_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03775_ VGND
+ VGND VPWR VPWR _03776_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12204_ _05139_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND
+ VGND VPWR VPWR _05289_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13184_ _06133_ _06135_ _06137_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__a21oi_2
X_10396_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _03711_ VGND
+ VGND VPWR VPWR _03713_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12135_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05225_ VGND
+ VGND VPWR VPWR _05226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12066_ _05165_ _05166_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a21oi_1
X_11017_ _04242_ _04246_ _04257_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12968_ _05939_ _05940_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__o21ai_2
X_14707_ clknet_leaf_51_i_clk net192 VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11919_ _05044_ _05040_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _05887_
+ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__xnor2_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14638_ clknet_leaf_59_i_clk _00183_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14569_ clknet_leaf_34_i_clk _00115_ VGND VGND VPWR VPWR diff2\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08090_ _01562_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08992_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _02476_
+ _02477_ _02414_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07943_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__buf_2
X_07874_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] _01488_ _01490_ _01453_
+ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__a31o_1
X_09613_ _03025_ _03022_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__o21bai_2
X_09544_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _02966_ VGND
+ VGND VPWR VPWR _02968_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09475_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02904_ VGND
+ VGND VPWR VPWR _02905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08426_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\] _01972_ VGND VGND VPWR
+ VPWR _01974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08357_ _01909_ _01910_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07308_ _01053_ _01054_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__and2_1
X_08288_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[17\] _01464_ VGND VGND VPWR
+ VPWR _01860_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07239_ _00998_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10250_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03572_ VGND
+ VGND VPWR VPWR _03595_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10181_ _03531_ _03532_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__nor2_1
X_13940_ _06431_ _06785_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__and2_1
X_13871_ _06725_ _06726_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _06554_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__a2bb2o_1
X_12822_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05789_ VGND
+ VGND VPWR VPWR _05826_ sky130_fd_sc_hd__xor2_2
XFILLER_0_97_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _05652_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04851_ VGND
+ VGND VPWR VPWR _04852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14423_ _07192_ _07199_ _07200_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__a21oi_1
X_11635_ _04773_ net476 _04792_ _04793_ _04788_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14354_ _01253_ _07141_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__and2_1
X_11566_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04723_ VGND
+ VGND VPWR VPWR _04740_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13305_ _06236_ _06237_ _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__a21oi_1
X_10517_ _03605_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03821_
+ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14285_ _07078_ _07081_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11497_ _04631_ _04651_ _04652_ _04666_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__or4_2
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13236_ _06176_ _06178_ _06181_ _05860_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__a31o_1
X_10448_ net117 _03719_ _03744_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13167_ _06122_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10379_ _03535_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__and2_1
X_12118_ _05206_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__xor2_1
X_13098_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__and2_1
X_12049_ _05139_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__clkbuf_4
X_07590_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[4\] _01277_ _01255_ VGND
+ VGND VPWR VPWR _01278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09260_ _02694_ _02718_ _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_157_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08211_ _01793_ _01795_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__nor2_1
X_09191_ _02649_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08142_ _01556_ _01727_ _01732_ _01733_ _01485_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08073_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08975_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _02461_ VGND
+ VGND VPWR VPWR _02462_ sky130_fd_sc_hd__xnor2_1
Xhold15 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND VGND
+ VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 _00710_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _01533_ _01535_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\]
+ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__a21oi_1
Xhold48 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND VPWR VPWR
+ net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[3\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[4\] VGND VGND VPWR VPWR _01477_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07788_ net18 _01423_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09527_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _02951_ VGND
+ VGND VPWR VPWR _02952_ sky130_fd_sc_hd__xor2_2
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09458_ _02888_ _02889_ _02755_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08409_ _01873_ _01959_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09389_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _02806_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__a311o_1
XFILLER_0_108_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11420_ _04442_ _04607_ _04608_ _04456_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11351_ _04547_ _04548_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10302_ _03280_ _03628_ _03629_ _03631_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14070_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06565_ _06899_
+ _06900_ _06631_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__o221a_1
X_11282_ _04484_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__or2_1
X_13021_ _05992_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10233_ _03575_ _03578_ _03580_ _03191_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10164_ _03499_ _03502_ _03511_ _03516_ _03510_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__o32a_1
X_14972_ clknet_leaf_89_i_clk _00517_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10095_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ _03205_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13923_ _06770_ _06771_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__xnor2_1
X_13854_ _06710_ _06711_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__nand2_1
X_12805_ _05632_ _05810_ _05811_ _05675_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13785_ _06650_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _06651_ sky130_fd_sc_hd__nor2_1
X_10997_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _04240_ VGND
+ VGND VPWR VPWR _04241_ sky130_fd_sc_hd__xnor2_1
X_12736_ _05737_ _05740_ _05748_ _05490_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__o31ai_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12667_ _05687_ _05688_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14406_ _01253_ _07186_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__and2_1
X_11618_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND VPWR
+ VPWR _04779_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15386_ clknet_leaf_47_i_clk _00931_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_12598_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _05626_ VGND
+ VGND VPWR VPWR _05628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14337_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _07125_ VGND
+ VGND VPWR VPWR _07126_ sky130_fd_sc_hd__xnor2_1
X_11549_ _04378_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND
+ VGND VPWR VPWR _04726_ sky130_fd_sc_hd__or2_1
Xhold507 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14268_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _07041_ VGND
+ VGND VPWR VPWR _07067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13219_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06136_ VGND
+ VGND VPWR VPWR _06168_ sky130_fd_sc_hd__xor2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14199_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _06646_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__o21ba_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _02270_ _02272_ _02277_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a21o_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ net9 _01366_ net10 VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__o21ai_1
X_08691_ _02199_ _02202_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__nand2_1
X_07642_ _01319_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07573_ _01264_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09312_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND VPWR
+ VPWR _02764_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09243_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _02704_ VGND
+ VGND VPWR VPWR _02705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09174_ _02641_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08125_ _01457_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _01651_ _01652_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08958_ _02445_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__nor2_1
X_07909_ _01328_ _01520_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__or2_1
X_08889_ _02319_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__clkbuf_4
X_10920_ _04155_ _04170_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__or2b_1
X_10851_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04109_ VGND
+ VGND VPWR VPWR _04110_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _06201_ _06468_ _06469_ _06459_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__o211a_1
X_10782_ _03669_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05556_
+ _05526_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__o21a_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ clknet_leaf_12_i_clk _00785_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _05500_ net350 _05495_ _05502_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11403_ _04593_ _04589_ _04590_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15171_ clknet_leaf_113_i_clk _00716_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_62_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12383_ _05142_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05446_
+ _05447_ _05391_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14122_ _06940_ _06942_ _06934_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__mux2_1
X_11334_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04518_ _04414_
+ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14053_ _06877_ _06884_ _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__a21oi_1
X_11265_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04469_ VGND
+ VGND VPWR VPWR _04470_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_76_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13004_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND
+ VPWR VPWR _05978_ sky130_fd_sc_hd__inv_2
X_10216_ _03563_ _03554_ _03556_ _03557_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__nand4_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11196_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04409_
+ _04391_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__o21ai_1
X_10147_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__inv_2
X_14955_ clknet_leaf_90_i_clk _00500_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10078_ _03024_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13906_ _06755_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__xnor2_1
X_14886_ clknet_leaf_108_i_clk _00431_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13837_ _06691_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_14_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13768_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _06625_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12719_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__or4_2
XFILLER_0_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13699_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _06576_
+ _06577_ _06569_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15438_ clknet_leaf_31_i_clk _00983_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_29_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15369_ clknet_leaf_29_i_clk _00914_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold304 net68 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold337 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[16\] VGND VGND VPWR VPWR
+ net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _03305_ VGND
+ VGND VPWR VPWR _03306_ sky130_fd_sc_hd__and2_1
Xhold359 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _03246_
+ _03183_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__a21o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _02319_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__buf_4
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _03186_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__clkbuf_4
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\] _02261_ VGND VGND VPWR
+ VPWR _02262_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _02002_ _02193_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ r_i_alpha1\[11\] _01305_ _01276_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__mux2_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07556_ _01251_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07487_ _01080_ _01119_ _01120_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09226_ _02322_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02687_
+ _02688_ _02689_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09157_ _02611_ _02620_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08108_ _01663_ _01701_ _01680_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09088_ _02563_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08039_ net37 net55 VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__or2b_2
X_11050_ _04023_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04288_
+ _04289_ _04059_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__o221a_1
XFILLER_0_101_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10001_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _03356_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__or3_2
X_14740_ clknet_leaf_65_i_clk _00285_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_11952_ _05074_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__and2b_1
X_10903_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14671_ clknet_leaf_55_i_clk _00216_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_11883_ _05012_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__clkbuf_1
X_13622_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06514_ VGND
+ VGND VPWR VPWR _06515_ sky130_fd_sc_hd__nand2_1
X_10834_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04094_ VGND
+ VGND VPWR VPWR _04095_ sky130_fd_sc_hd__xor2_2
XFILLER_0_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13553_ _06451_ _06453_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10765_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ _05203_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05535_ _05545_
+ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__o41a_1
XFILLER_0_109_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13484_ _06392_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__nor2_1
X_10696_ _03981_ _03982_ _03983_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15223_ clknet_leaf_16_i_clk _00768_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12435_ _05488_ net237 _05141_ _05491_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15154_ clknet_leaf_115_i_clk _00699_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12366_ _05431_ _05432_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__or2b_1
X_14105_ _06909_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__clkbuf_4
X_11317_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15085_ clknet_leaf_119_i_clk _00630_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_12297_ _05363_ _05357_ _05368_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__a21oi_1
X_14036_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06837_ VGND
+ VGND VPWR VPWR _06871_ sky130_fd_sc_hd__nand2_1
X_11248_ _01251_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11179_ _04061_ _04393_ _04394_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14938_ clknet_leaf_109_i_clk net187 VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14869_ clknet_leaf_84_i_clk _00414_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_07410_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ _01132_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__or3_1
X_08390_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[14\] _01942_ _01943_
+ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07341_ _01056_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07272_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR _01021_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09011_ _02486_ _02490_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold112 net83 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold145 diff2\[15\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net107 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _03291_ sky130_fd_sc_hd__or2_1
Xhold178 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 net102 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _03226_
+ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _03168_ _03176_ _02132_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08726_ _02241_ _02235_ _02246_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__a21oi_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\] _02182_ VGND VGND VPWR
+ VPWR _02184_ sky130_fd_sc_hd__or2_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07608_ _01273_ diff1\[8\] VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__and2_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[16\] _02111_ VGND VGND VPWR
+ VPWR _02122_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07539_ net375 net236 _01234_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ _03848_ _03850_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09209_ _02237_ _02673_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__or2_1
X_10481_ _03789_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12220_ _05295_ _05299_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12151_ _05239_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11102_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04325_ VGND
+ VGND VPWR VPWR _04337_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12082_ _05130_ _05180_ _05181_ _05080_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__o211a_1
X_11033_ _04258_ _04273_ _04265_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__o21bai_2
X_12984_ _05952_ _05959_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11935_ _04795_ _05059_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14723_ clknet_leaf_55_i_clk _00268_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14654_ clknet_leaf_49_i_clk _00199_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _04757_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__nor2_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13605_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06499_
+ _06500_ _06285_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__o221a_1
X_10817_ _04072_ _04073_ _04078_ _03996_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14585_ clknet_leaf_35_i_clk _00130_ VGND VGND VPWR VPWR diff3\[10\] sky130_fd_sc_hd__dfxtp_1
X_11797_ _04557_ _04915_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13536_ _06437_ _06438_ _06205_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__o21ai_1
X_10748_ _04016_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13467_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _06351_ VGND
+ VGND VPWR VPWR _06379_ sky130_fd_sc_hd__xnor2_1
X_10679_ _03967_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15206_ clknet_leaf_1_i_clk _00751_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12418_ _05474_ _05476_ _01249_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__o21a_1
X_13398_ _06316_ _06317_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15137_ clknet_leaf_125_i_clk _00682_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12349_ _05378_ _05388_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15068_ clknet_leaf_102_i_clk _00613_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14019_ _06856_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
X_07890_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\] _01504_ _01464_ VGND
+ VGND VPWR VPWR _01505_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09560_ _02969_ _02975_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08511_ _02050_ _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__nor2_1
X_09491_ _02771_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08442_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _01988_ _01868_
+ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08373_ _01926_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07324_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _01038_ VGND VGND
+ VPWR VPWR _01069_ sky130_fd_sc_hd__or4_4
XFILLER_0_34_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07255_ _01007_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09827_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _03218_
+ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__xnor2_1
X_09758_ _03161_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\]
+ _02208_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__or3_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03097_ VGND
+ VGND VPWR VPWR _03098_ sky130_fd_sc_hd__xor2_2
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _04865_ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__or2_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _04802_
+ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__or2_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10602_ _03882_ _03891_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14370_ _07143_ _07139_ _07147_ _07152_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11582_ _04753_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13321_ _06202_ _06250_ _06252_ _06110_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10533_ _03623_ _03834_ _03835_ _03780_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13252_ _04538_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10464_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03774_ VGND
+ VGND VPWR VPWR _03775_ sky130_fd_sc_hd__xor2_2
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12203_ _05285_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06136_ VGND
+ VGND VPWR VPWR _06137_ sky130_fd_sc_hd__xnor2_1
X_10395_ _03711_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _03712_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05163_ VGND VGND VPWR
+ VPWR _05225_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12065_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR _05167_ sky130_fd_sc_hd__inv_2
X_11016_ _04258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12967_ _05943_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11918_ _05038_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__inv_2
X_14706_ clknet_leaf_50_i_clk net156 VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12898_ _05884_ _05886_ _05878_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__mux2_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11849_ _04980_ _04981_ _04786_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__o21ai_1
X_14637_ clknet_leaf_43_i_clk _00182_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14568_ clknet_leaf_34_i_clk _00114_ VGND VGND VPWR VPWR diff2\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13519_ _06210_ net330 _06203_ _06423_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__o211a_1
X_14499_ clknet_leaf_4_i_clk _00045_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08991_ _02463_ _02466_ _02475_ _02369_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__a31o_1
X_07942_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _01549_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07873_ _01488_ _01490_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] VGND
+ VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a21oi_1
X_09612_ _02591_ _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09543_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _02966_ VGND
+ VGND VPWR VPWR _02967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09474_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _02903_ VGND
+ VGND VPWR VPWR _02904_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08425_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\] _01972_ VGND VGND VPWR
+ VPWR _01973_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08356_ _01550_ _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07307_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _01038_ VGND
+ VGND VPWR VPWR _01054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08287_ _01857_ _01858_ _01562_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07238_ net368 net19 _00993_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10180_ _03519_ _03526_ _03524_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__o21ai_1
X_13870_ _06722_ _06721_ _06723_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__o21ba_1
X_12821_ _05825_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12752_ _05486_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _05762_
+ _05764_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__a22o_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _04794_ VGND VGND VPWR
+ VPWR _04851_ sky130_fd_sc_hd__o31a_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05501_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _05701_
+ _05702_ _05544_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__o221a_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _07144_ VGND
+ VGND VPWR VPWR _07200_ sky130_fd_sc_hd__xor2_1
X_11634_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _04791_
+ _04786_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14353_ _06903_ _07138_ _07139_ _07140_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__o31ai_1
X_11565_ _04376_ _04737_ _04738_ _04739_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13304_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR _06238_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10516_ _03817_ _03820_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14284_ _07057_ _07079_ _07080_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11496_ _04651_ _04655_ _04666_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13235_ _06176_ _06178_ _06181_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__a21oi_1
X_10447_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13166_ _06069_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__and2_1
X_10378_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _03696_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__mux2_1
X_12117_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _05209_ VGND
+ VGND VPWR VPWR _05210_ sky130_fd_sc_hd__xnor2_1
X_13097_ _05998_ _06058_ _06059_ _05938_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12048_ _05140_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _05151_ _05152_ _04965_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__o221a_1
X_13999_ _06834_ _06836_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08210_ _01529_ net542 _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__o21ai_1
X_09190_ _02655_ _02656_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08141_ _01722_ _01731_ _01572_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08072_ _01662_ _01663_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08974_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ _02442_ _02342_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__o31a_1
Xhold16 _00423_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 _00593_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] _01534_ VGND VGND
+ VPWR VPWR _01535_ sky130_fd_sc_hd__nand2_1
Xhold38 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[3\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[4\] VGND VGND VPWR VPWR _01476_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07787_ _01423_ _01424_ net247 _01333_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__o2bb2a_1
X_09526_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _02771_ _02937_
+ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09457_ _02874_ _02881_ _02887_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__nor3_1
XFILLER_0_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08408_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__buf_2
X_09388_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02813_
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08339_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] _01900_ _01869_
+ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11350_ _04540_ _04546_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10301_ _03605_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11281_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04483_ VGND
+ VGND VPWR VPWR _04485_ sky130_fd_sc_hd__nor2_1
X_13020_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _05982_ VGND
+ VGND VPWR VPWR _05993_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10232_ _03561_ _03564_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a21o_1
X_10163_ _03497_ _03509_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__nor2_1
X_14971_ clknet_leaf_105_i_clk _00516_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10094_ _03389_ _03452_ _03453_ _03292_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__o211a_1
X_13922_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _06716_ VGND
+ VGND VPWR VPWR _06771_ sky130_fd_sc_hd__xnor2_1
X_13853_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _06707_ _06694_
+ _06698_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__a211oi_1
X_12804_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _05811_ sky130_fd_sc_hd__or2_1
X_10996_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04034_ VGND VGND VPWR
+ VPWR _04240_ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13784_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND
+ VPWR VPWR _06650_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12735_ _05737_ _05740_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__o21a_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _05641_ VGND
+ VGND VPWR VPWR _05688_ sky130_fd_sc_hd__xor2_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND VPWR
+ VPWR _04778_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14405_ _06903_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _07184_
+ _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__a22o_1
X_12597_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _05626_ VGND
+ VGND VPWR VPWR _05627_ sky130_fd_sc_hd__and2_1
X_15385_ clknet_leaf_29_i_clk _00930_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11548_ _04722_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14336_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _07125_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_135_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold508 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14267_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _07042_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__o21ai_1
Xhold519 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR
+ VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11479_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04661_ VGND
+ VGND VPWR VPWR _04662_ sky130_fd_sc_hd__xor2_1
X_13218_ _05998_ _06166_ _06167_ _06110_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14198_ _06905_ _07004_ _07005_ _06996_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__o211a_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _06096_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _06106_ sky130_fd_sc_hd__and2b_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ net9 net10 _01366_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__or3_1
X_08690_ _02161_ _02165_ _02176_ _02185_ _02204_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__o2111a_1
X_07641_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\] _01318_ _01282_
+ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__mux2_1
X_07572_ net250 net450 _01255_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__mux2_1
X_09311_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND VPWR
+ VPWR _02763_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09242_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _02703_ VGND
+ VGND VPWR VPWR _02704_ sky130_fd_sc_hd__xor2_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09173_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _02640_ VGND
+ VGND VPWR VPWR _02641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08124_ _01539_ net596 _01713_ _01716_ _01661_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08055_ net38 net56 VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08957_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _02444_ VGND
+ VGND VPWR VPWR _02446_ sky130_fd_sc_hd__nor2_1
X_07908_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[11\]
+ _01508_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__and3_1
X_08888_ _02321_ net447 _02381_ _02386_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07839_ net164 _01457_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__or2_1
X_10850_ _04034_ _04108_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _02921_ _02930_ _02934_ _02761_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__a31o_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04042_
+ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12520_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _05558_ _05559_ _05544_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _05501_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11402_ _04589_ _04590_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__o21ai_1
X_15170_ clknet_leaf_113_i_clk _00715_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12382_ _05438_ _05441_ _05445_ _05222_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14121_ _06941_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__inv_2
X_11333_ _04442_ _04531_ _04532_ _04456_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14052_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06845_ VGND
+ VGND VPWR VPWR _06885_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11264_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04412_ VGND VGND VPWR
+ VPWR _04469_ sky130_fd_sc_hd__o31a_1
X_13003_ _05871_ net411 _05976_ _05977_ _05910_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__o221a_1
X_10215_ _03554_ _03556_ _03557_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11195_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04409_
+ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__and2_1
X_10146_ _03480_ _03487_ _03489_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a21oi_1
X_14954_ clknet_leaf_89_i_clk _00499_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10077_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03439_ _03185_
+ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__mux2_1
X_13905_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06716_ _06752_
+ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__a21o_1
X_14885_ clknet_leaf_110_i_clk net125 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13836_ _06694_ _06695_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10979_ _04223_ _04224_ _04012_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__o21ai_1
X_13767_ _06556_ _06635_ _06636_ _06459_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12718_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _05733_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13698_ _06576_ _06577_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15437_ clknet_leaf_27_i_clk _00982_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_12649_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _05674_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15368_ clknet_leaf_21_i_clk _00913_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_142_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold305 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ _07109_ _07110_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold316 _01247_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ clknet_leaf_17_i_clk _00844_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold327 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold338 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 diff1\[17\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09860_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _03246_
+ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__nor2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _02320_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__clkbuf_4
X_09791_ _03184_ net226 _03017_ _03188_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__o211a_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\] _02249_ _01881_ VGND
+ VGND VPWR VPWR _02261_ sky130_fd_sc_hd__o21a_1
X_08673_ _02198_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
X_07624_ diff2\[11\] _01270_ _01272_ diff3\[11\] _01304_ VGND VGND VPWR VPWR _01305_
+ sky130_fd_sc_hd__a221o_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ net1 VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07486_ _01016_ net253 _01207_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09225_ _02308_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__buf_4
XFILLER_0_29_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09156_ _02322_ net548 _02623_ _02625_ _02414_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08107_ _01679_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__inv_2
X_09087_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _02555_ VGND
+ VGND VPWR VPWR _02564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08038_ net55 net37 VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__or2b_2
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10000_ _03237_ net550 _03368_ _03369_ _03258_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__o221a_1
X_09989_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03358_ VGND
+ VGND VPWR VPWR _03360_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11951_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05072_ _05073_
+ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10902_ _04142_ _04144_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a21oi_1
X_11882_ _05011_ _03118_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__and2b_1
X_14670_ clknet_leaf_54_i_clk _00215_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10833_ _04034_ _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__nand2_1
X_13621_ _06488_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10764_ _04033_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__buf_2
X_13552_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06452_ VGND
+ VGND VPWR VPWR _06453_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _05203_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _05539_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__nand3_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13483_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06337_ VGND
+ VGND VPWR VPWR _06393_ sky130_fd_sc_hd__xnor2_1
X_10695_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _03944_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12434_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _05490_
+ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__or2_1
X_15222_ clknet_leaf_16_i_clk _00767_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15153_ clknet_leaf_123_i_clk _00698_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_12365_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05430_ VGND
+ VGND VPWR VPWR _05432_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11316_ _04431_ net544 _04515_ _04516_ _04360_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14104_ _06910_ net303 _06925_ _06927_ _06922_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__o221a_1
X_15084_ clknet_leaf_120_i_clk _00629_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_12296_ _05363_ _05357_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14035_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06837_ VGND
+ VGND VPWR VPWR _06870_ sky130_fd_sc_hd__or2_1
X_11247_ _04444_ net583 VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__or2_1
X_11178_ _04375_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__buf_4
X_10129_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03477_ _03205_
+ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__o21a_1
X_14937_ clknet_leaf_110_i_clk _00482_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14868_ clknet_leaf_84_i_clk _00413_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06680_ VGND
+ VGND VPWR VPWR _06681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14799_ clknet_leaf_72_i_clk _00344_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07340_ _01082_ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07271_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09010_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _02493_ VGND
+ VGND VPWR VPWR _02494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold102 _00651_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 net96 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _00480_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net252 sky130_fd_sc_hd__buf_1
XFILLER_0_110_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold146 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09912_ _03185_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__buf_2
Xhold179 _00823_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _03228_
+ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__nand2_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _03174_ _03175_ _02804_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_60_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08725_ _02244_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__nor2_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\] _02182_ VGND VGND VPWR
+ VPWR _02183_ sky130_fd_sc_hd__and2_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07607_ _01291_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _02103_ _02106_ _02114_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__nand3_1
XFILLER_0_95_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_75_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07538_ _01241_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07469_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _01045_ _01088_
+ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _02672_ VGND
+ VGND VPWR VPWR _02673_ sky130_fd_sc_hd__xor2_1
X_10480_ _03787_ _03788_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09139_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02609_ VGND
+ VGND VPWR VPWR _02610_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12150_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _05238_ VGND
+ VGND VPWR VPWR _05240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11101_ _04310_ _04332_ _04333_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_13_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12081_ _05132_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11032_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _04263_ _04254_
+ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_28_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12983_ _05944_ _05946_ _05954_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__a21bo_1
X_14722_ clknet_leaf_53_i_clk _00267_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_11934_ _04970_ _05025_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ clknet_leaf_49_i_clk net308 VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _04996_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _06490_ _06495_ _06498_ _06216_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__a31o_1
X_10816_ _04072_ _04073_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__o21ai_1
X_11796_ _04557_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04915_
+ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14584_ clknet_leaf_36_i_clk _00129_ VGND VGND VPWR VPWR diff3\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13535_ _06421_ _06428_ _06427_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10747_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10678_ _03954_ _03962_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__nand2_1
X_13466_ _06372_ _06378_ _01766_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_153_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15205_ clknet_leaf_1_i_clk _00750_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12417_ _05474_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13397_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _06315_ VGND
+ VGND VPWR VPWR _06317_ sky130_fd_sc_hd__or2_1
X_15136_ clknet_leaf_122_i_clk _00681_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_12348_ _05397_ _05414_ _05409_ _05415_ _05408_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__o32a_1
X_15067_ clknet_leaf_117_i_clk _00612_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_12279_ _05348_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _05353_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14018_ _01253_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08510_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\] _02049_ VGND VGND VPWR
+ VPWR _02051_ sky130_fd_sc_hd__and2b_1
X_09490_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ _02882_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__or4_2
XFILLER_0_81_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08441_ _01986_ _01987_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08372_ _01927_ _01928_ _01882_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07323_ _01047_ _01066_ _01067_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07254_ net386 net9 _01000_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09826_ _02851_ _03216_ _03217_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__a21bo_1
X_09757_ _03024_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__and2_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _02213_ _02223_ _02222_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__or3_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03087_ _02770_
+ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__o21a_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08639_ _02167_ _01979_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__and2b_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _04769_ net560 _04762_ _04806_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__o211a_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10601_ _03865_ _03872_ _03877_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__a21o_1
X_11581_ _04391_ _02310_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10532_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _03835_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13320_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13251_ _06185_ _06193_ _06194_ _05860_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__a31o_1
X_10463_ _03651_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12202_ _05286_ _05282_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__or2b_1
X_13182_ _06112_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__clkbuf_4
X_10394_ _03708_ _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12133_ _05224_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12064_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _05148_ _05164_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a31o_1
X_11015_ _04242_ _04246_ _04257_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12966_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05942_ VGND
+ VGND VPWR VPWR _05944_ sky130_fd_sc_hd__nand2_1
X_14705_ clknet_leaf_56_i_clk _00250_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_2
X_11917_ _05043_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__inv_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ clknet_leaf_43_i_clk _00181_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14567_ clknet_leaf_35_i_clk _00113_ VGND VGND VPWR VPWR diff2\[11\] sky130_fd_sc_hd__dfxtp_1
X_11779_ _04907_ _04910_ _04919_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13518_ _06421_ _06422_ _06232_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__o21ai_1
X_14498_ clknet_leaf_25_i_clk _00044_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13449_ _06362_ _06363_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15119_ clknet_leaf_116_i_clk _00664_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_08990_ _02463_ _02466_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__a21oi_1
X_07941_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[16\] _01544_ _01543_
+ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07872_ _01328_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__nand2_1
X_09611_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _03026_ VGND
+ VGND VPWR VPWR _03027_ sky130_fd_sc_hd__xnor2_1
X_09542_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _02965_ VGND
+ VGND VPWR VPWR _02966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09473_ _02770_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08424_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[3\] _01971_ VGND VGND VPWR
+ VPWR _01972_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08355_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] _01898_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND VPWR VPWR _01914_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07306_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _01038_ VGND
+ VGND VPWR VPWR _01053_ sky130_fd_sc_hd__or2_1
X_08286_ _01746_ _01852_ _01770_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07237_ _00997_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09809_ _03198_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__inv_2
X_12820_ _05652_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _05485_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nor2_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _01252_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__buf_2
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12682_ _05694_ _05696_ _05700_ _05486_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__a31o_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _07196_ _07193_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__or2b_1
X_11633_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _04791_
+ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__and2_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14352_ _06903_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND
+ VGND VPWR VPWR _07140_ sky130_fd_sc_hd__nand2_1
X_11564_ _04455_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_887 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13303_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _06218_ _06235_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__a31o_1
X_10515_ _03817_ _03820_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__nand2_1
X_11495_ _04649_ _04663_ _04664_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__a21o_1
X_14283_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _07041_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__o41ai_4
XFILLER_0_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13234_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06142_ VGND
+ VGND VPWR VPWR _06181_ sky130_fd_sc_hd__xor2_1
X_10446_ _03626_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _03757_
+ _03758_ _03633_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13165_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06120_ _05844_
+ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__mux2_1
X_10377_ _03694_ _03695_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12116_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05208_ VGND
+ VGND VPWR VPWR _05209_ sky130_fd_sc_hd__xnor2_1
X_13096_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _06059_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12047_ _05146_ _05150_ _05129_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13998_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06837_ VGND
+ VGND VPWR VPWR _06838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12949_ _05843_ _05926_ _05929_ _05675_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14619_ clknet_leaf_44_i_clk _00164_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08140_ _01722_ _01731_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08071_ _01664_ _01666_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08973_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02458_ _02459_
+ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold17 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[13\]
+ _01520_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__or3_1
Xhold39 _00251_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\] _01471_
+ _01473_ _01475_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__o221a_1
X_07786_ net17 _01421_ _01344_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09525_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02938_ VGND
+ VGND VPWR VPWR _02950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09456_ _02874_ _02881_ _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08407_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR _02828_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08338_ _01550_ _01897_ _01899_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08269_ _01529_ net551 _01794_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10300_ _03628_ _03629_ _03280_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11280_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04483_ VGND
+ VGND VPWR VPWR _04484_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10231_ _03574_ _03576_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10162_ _03389_ _03513_ _03514_ _03515_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__o211a_1
X_14970_ clknet_leaf_105_i_clk _00515_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_10093_ _03290_ net620 VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__or2_1
X_13921_ _06761_ _06766_ _06760_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ _06671_ _06679_ _06687_ _06691_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ _05806_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__xor2_1
X_13783_ _06561_ _06647_ _06485_ _06649_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__o211a_1
X_10995_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _04239_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _05746_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12665_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05648_ _05684_
+ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14404_ _07183_ _07179_ _07180_ _01861_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__o31a_1
X_11616_ _04773_ net509 _04776_ _04777_ _04539_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__o221a_1
X_15384_ clknet_leaf_47_i_clk _00929_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12596_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05625_ VGND
+ VGND VPWR VPWR _05626_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14335_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _07124_ sky130_fd_sc_hd__inv_2
X_11547_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04723_ _04719_
+ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold509 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _07042_ _07057_
+ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__o21bai_1
X_11478_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] net652 _04412_ VGND
+ VGND VPWR VPWR _04661_ sky130_fd_sc_hd__o41a_1
XFILLER_0_111_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13217_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _06167_ sky130_fd_sc_hd__or2_1
X_10429_ _03741_ _03742_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14197_ _06907_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _07005_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _06103_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nor2_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06003_ VGND
+ VGND VPWR VPWR _06044_ sky130_fd_sc_hd__xnor2_1
X_07640_ r_i_alpha1\[14\] _01317_ _01258_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07571_ _01263_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09310_ _02757_ net280 _02760_ _02762_ _02689_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09241_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02695_ _02343_
+ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09172_ _02498_ _02639_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08123_ _01472_ _01715_ _01480_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ net56 net38 VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08956_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _02444_ VGND
+ VGND VPWR VPWR _02445_ sky130_fd_sc_hd__and2_1
X_07907_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[11\] _01518_
+ _01519_ _01513_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__o221a_1
X_08887_ _02382_ _02384_ _02385_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _02320_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__o221ai_1
X_07838_ _01454_ net250 _01460_ _01461_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07769_ _01273_ _01413_ _01411_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__mux2_1
X_09508_ _02921_ _02930_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__a21oi_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10780_ _04047_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__clkbuf_4
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _02769_ VGND VGND VPWR
+ VPWR _02872_ sky130_fd_sc_hd__o31a_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _05489_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11401_ _04591_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12381_ _05438_ _05441_ _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14120_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _06929_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__or3_1
X_11332_ _04444_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _04532_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14051_ _06878_ _06880_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11263_ _01252_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13002_ _05973_ _05975_ _05845_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__o21ai_1
X_10214_ _03561_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__nand2_1
X_11194_ _04407_ _04408_ _04061_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__mux2_1
X_10145_ _03482_ _03488_ _03489_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14953_ clknet_leaf_104_i_clk _00498_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10076_ _03433_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13904_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06707_ VGND
+ VGND VPWR VPWR _06755_ sky130_fd_sc_hd__xnor2_1
X_14884_ clknet_leaf_110_i_clk net127 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13835_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _06684_ VGND
+ VGND VPWR VPWR _06695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13766_ _06557_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__or2_1
X_10978_ _04216_ _04222_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12717_ _05725_ _05728_ _05724_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__a21oi_2
X_13697_ _06292_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _06567_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15436_ clknet_leaf_27_i_clk _00981_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_12648_ _05671_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15367_ clknet_leaf_21_i_clk _00912_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_12579_ _05597_ _05603_ _05601_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14318_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _07042_ VGND
+ VGND VPWR VPWR _07110_ sky130_fd_sc_hd__xnor2_1
X_15298_ clknet_leaf_14_i_clk _00843_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold306 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 net72 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold328 diff2\[4\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold339 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14249_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _07023_ VGND
+ VGND VPWR VPWR _07051_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__clkbuf_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ net132 _03186_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__or2_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _01866_ _02258_ _02259_ _02260_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__o211a_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _01981_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__and2_1
X_07623_ _01273_ diff1\[11\] VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__and2_1
X_07554_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07485_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _01159_ _01205_
+ _01206_ _01030_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09224_ _02674_ _02682_ _02686_ _02313_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09155_ _02320_ _02624_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08106_ _01664_ _01681_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__nand2_2
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09086_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _02555_ VGND
+ VGND VPWR VPWR _02563_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08037_ _01455_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09988_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03358_ VGND
+ VGND VPWR VPWR _03359_ sky130_fd_sc_hd__nand2_1
X_08939_ _02429_ _01979_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__and2b_1
X_11950_ _05072_ _05073_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ _04142_ _04144_ _04135_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__o21a_1
X_11881_ _04770_ _05000_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__o21a_1
X_13620_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06488_ VGND
+ VGND VPWR VPWR _06513_ sky130_fd_sc_hd__or2_1
X_10832_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__or4_1
X_13551_ _06234_ _06410_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__nand2_1
X_10763_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _04033_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12502_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _05542_ _05543_ _05544_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13482_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06352_ _06389_
+ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__a21o_1
X_10694_ _03960_ _03961_ _03980_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15221_ clknet_leaf_16_i_clk _00766_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12433_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15152_ clknet_leaf_123_i_clk _00697_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12364_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _05430_ VGND
+ VGND VPWR VPWR _05431_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14103_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _06923_
+ _06924_ _06926_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__a31o_1
X_11315_ _04503_ _04506_ _04514_ _04396_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__a31o_1
X_15083_ clknet_leaf_99_i_clk _00628_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _05366_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14034_ _06866_ _06863_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__or2b_1
X_11246_ _04448_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__xor2_1
X_11177_ _04393_ _04394_ _04061_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__a21oi_2
X_10128_ _03389_ _03483_ _03484_ _03292_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14936_ clknet_leaf_110_i_clk _00481_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10059_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03423_ _03185_
+ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__mux2_1
X_14867_ clknet_leaf_84_i_clk _00412_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13818_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__nor4_1
X_14798_ clknet_leaf_71_i_clk _00343_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13749_ _06292_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _06615_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07270_ _01018_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15419_ clknet_leaf_24_i_clk _00964_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold103 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold114 net80 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold125 CORDIC_PE\[0\].genblk1.cordic_engine_inst.i_quadrant\[1\] VGND VGND VPWR
+ VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold136 net77 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold158 _00601_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _03284_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__xor2_1
Xhold169 _00545_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ net298 _03189_ _03230_ _03231_ _03013_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__o221a_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _03173_ _03170_ _03171_ _03172_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__or4_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_9_i_clk sky130_fd_sc_hd__clkbuf_16
X_08724_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\] _02243_ VGND VGND VPWR
+ VPWR _02245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\] _02181_ VGND VGND VPWR
+ VPWR _02182_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[7\] _01290_ _01282_ VGND
+ VGND VPWR VPWR _01291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\] _02113_ _02119_ VGND
+ VGND VPWR VPWR _02120_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07537_ net372 net322 _01234_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07468_ _01076_ _01084_ _01079_ _01080_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09207_ _02343_ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07399_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09138_ _02342_ _02608_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09069_ _02542_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__nand2_1
X_11100_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04316_ _04327_
+ _04334_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a31o_1
X_12080_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05179_
+ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__xor2_1
X_11031_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _04271_ VGND
+ VGND VPWR VPWR _04272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12982_ _05958_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
X_14721_ clknet_leaf_53_i_clk _00266_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11933_ _05005_ _05009_ _05044_ _05057_ _05052_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__o2111ai_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ clknet_leaf_48_i_clk _00197_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _04989_ _04987_ _04993_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__or3b_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _06490_ _06495_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__a21oi_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _04076_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__and2_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ clknet_leaf_36_i_clk _00128_ VGND VGND VPWR VPWR diff3\[8\] sky130_fd_sc_hd__dfxtp_1
X_11795_ _04771_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04933_
+ _04934_ _04788_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13534_ _06435_ _06436_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__nor2_1
X_10746_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND VPWR
+ VPWR _04019_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13465_ _06200_ _06376_ _06377_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ _03965_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__nand2_1
X_15204_ clknet_leaf_1_i_clk _00749_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12416_ _05464_ _05461_ _05469_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13396_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _06315_ VGND
+ VGND VPWR VPWR _06316_ sky130_fd_sc_hd__and2_1
X_15135_ clknet_leaf_125_i_clk _00680_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12347_ _05395_ _05407_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15066_ clknet_leaf_117_i_clk net523 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12278_ _05140_ net321 _05141_ _05352_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__o211a_1
X_14017_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06854_ _06553_
+ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__mux2_1
X_11229_ _04437_ _04438_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14919_ clknet_leaf_87_i_clk _00464_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_08440_ _01974_ _01976_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08371_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[9\] _01914_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[10\]
+ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07322_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _01048_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07253_ _01006_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09825_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _03204_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _03217_ sky130_fd_sc_hd__a31o_1
X_09756_ _03158_ _03159_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _02746_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__a2bb2o_1
X_08707_ _02228_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__inv_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _02748_ _03095_ _03096_ _03058_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__o211a_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _01869_ _02156_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__o21a_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _02091_ _02094_ _02104_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10600_ _03606_ _03895_ _03896_ _03780_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11580_ _04376_ _04751_ _04752_ _04739_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10531_ _03828_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13250_ _06185_ _06193_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10462_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03760_ VGND
+ VGND VPWR VPWR _03773_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12201_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _05280_ VGND
+ VGND VPWR VPWR _05286_ sky130_fd_sc_hd__and2_1
X_13181_ _06085_ _06089_ _06117_ _06134_ _06131_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10393_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03709_ _03650_
+ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12132_ _04850_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12063_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _05158_
+ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__o21ai_1
X_11014_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12965_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05942_ VGND
+ VGND VPWR VPWR _05943_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11916_ _04850_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__and2_1
X_14704_ clknet_leaf_57_i_clk _00249_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12896_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _05872_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__or3_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ clknet_leaf_59_i_clk _00180_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__and2_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ clknet_leaf_35_i_clk _00112_ VGND VGND VPWR VPWR diff2\[10\] sky130_fd_sc_hd__dfxtp_1
X_11778_ _04907_ _04910_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13517_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10729_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _03999_
+ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14497_ clknet_leaf_4_i_clk _00043_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13448_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _06337_ VGND
+ VGND VPWR VPWR _06363_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13379_ _06296_ _06300_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__xor2_1
X_15118_ clknet_leaf_114_i_clk _00663_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15049_ clknet_leaf_111_i_clk net129 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_07940_ _01539_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[16\] _01546_
+ _01547_ _01513_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_74_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07871_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[4\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[5\]
+ _01469_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__or3_1
X_09610_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ _02769_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_89_i_clk clknet_4_5_0_i_clk VGND VGND VPWR VPWR clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09541_ _02771_ _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__and2_1
X_09472_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ _02882_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08423_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\]
+ _01549_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_12_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08354_ _01876_ net398 _01823_ _01913_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07305_ _01037_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08285_ _01746_ _01770_ _01852_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07236_ net341 net18 _00993_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09808_ net130 _03189_ _03200_ _03202_ _03013_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09739_ _03132_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__inv_2
X_12750_ _05732_ _05752_ _05754_ _05761_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__o211a_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _04849_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12681_ _05694_ _05696_ _05700_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__a21oi_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _07059_ _07197_ _07198_ _01475_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__o211a_1
X_11632_ _04789_ _04790_ _04445_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14351_ _07128_ _07130_ _07137_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11563_ _04378_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND
+ VGND VPWR VPWR _04738_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13302_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _06228_
+ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__o21ai_1
X_10514_ _03818_ _03819_ _03804_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__or3b_1
X_14282_ _07061_ _07067_ _07072_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11494_ _04674_ _04675_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__or2_2
XFILLER_0_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13233_ _06171_ _06180_ _01766_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10445_ _03755_ _03756_ _03631_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13164_ _06117_ _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__xnor2_1
X_10376_ _03683_ _03687_ _03684_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12115_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__and2b_1
X_13095_ _06056_ _06057_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12046_ _05146_ _05150_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13997_ _06807_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12948_ _05848_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12879_ _05854_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _05869_ _05870_ _05751_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__o221a_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14618_ clknet_leaf_44_i_clk _00163_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14549_ clknet_leaf_35_i_clk _00095_ VGND VGND VPWR VPWR diff1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08070_ _01653_ _01655_ _01665_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08972_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02458_ _02445_
+ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__a21o_1
X_07923_ _01532_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__inv_2
Xhold18 _00598_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _00365_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07854_ _01474_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07785_ net17 _01421_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__or2_1
X_09524_ _02949_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09455_ _02885_ _02886_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nor2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08406_ _01956_ _01953_ _01952_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_143_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09386_ _02757_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _02825_ _02826_ _02827_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08337_ _01550_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08268_ _01572_ _01727_ _01841_ _01842_ _01457_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08199_ _01563_ _01782_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__nor2_1
X_10230_ _03577_ _03564_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10161_ _01474_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__buf_4
X_10092_ _03446_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__xor2_1
X_13920_ _06769_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
X_13851_ _06696_ _06703_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12802_ _05807_ _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__or2_1
X_13782_ _06642_ _06648_ _06584_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__o21ai_2
X_10994_ _04227_ _04229_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12733_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _05745_ VGND
+ VGND VPWR VPWR _05747_ sky130_fd_sc_hd__or2_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05679_ _05686_ _04961_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__o21a_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14403_ _07179_ _07180_ _07183_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__o21ai_1
X_11615_ _04445_ _04774_ _04775_ _04755_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15383_ clknet_leaf_38_i_clk _00928_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12595_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05598_ _05525_ VGND
+ VGND VPWR VPWR _05625_ sky130_fd_sc_hd__o41a_1
X_14334_ _07117_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _07123_ sky130_fd_sc_hd__or2b_1
X_11546_ _04692_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14265_ _06905_ _07063_ _07064_ _06996_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__o211a_1
X_11477_ _04649_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__inv_2
X_13216_ _06164_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__and2_1
X_10428_ _03699_ _03724_ _03725_ _03734_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__nand4_2
X_14196_ _06999_ _07003_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__xor2_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _06100_ _06102_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__and2_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _03631_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] VGND
+ VGND VPWR VPWR _03679_ sky130_fd_sc_hd__and2_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _06043_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
X_12029_ _05130_ net205 _04979_ _05137_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07570_ net242 _01262_ _01255_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09240_ _02314_ _02701_ _02702_ _02260_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09171_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02608_ _02627_
+ _02342_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08122_ _01709_ _01714_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08053_ _01463_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[8\] _01635_ _01650_
+ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ _02441_ _02443_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__xnor2_1
X_07906_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[11\] _01517_ _01480_
+ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__a21o_1
X_08886_ _01959_ _02383_ _02382_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__a21oi_1
X_07837_ net165 _01457_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07768_ net11 _01408_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09507_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _02933_ VGND
+ VGND VPWR VPWR _02934_ sky130_fd_sc_hd__xnor2_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07699_ _01363_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09438_ _02871_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09369_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _02808_
+ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04565_ VGND
+ VGND VPWR VPWR _04592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12380_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05430_ VGND
+ VGND VPWR VPWR _05445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11331_ _04528_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14050_ _06883_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
X_11262_ _04467_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13001_ _05973_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__and2_1
X_10213_ _03558_ _03560_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__nand2_1
X_11193_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _04398_
+ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10144_ _03497_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14952_ clknet_leaf_106_i_clk _00497_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10075_ _03403_ _03435_ _03436_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__o211a_1
X_13903_ _06754_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
X_14883_ clknet_leaf_110_i_clk _00428_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13834_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _06684_ VGND
+ VGND VPWR VPWR _06694_ sky130_fd_sc_hd__and2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13765_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _06634_
+ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__xor2_1
X_10977_ _04216_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nor2_1
X_12716_ _05731_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
X_13696_ _06293_ _06571_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12647_ _05669_ _05670_ _05668_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15435_ clknet_leaf_27_i_clk _00980_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15366_ clknet_leaf_21_i_clk _00911_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12578_ _05608_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11529_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04694_ VGND
+ VGND VPWR VPWR _04708_ sky130_fd_sc_hd__nand2_1
X_14317_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _07042_ _07106_
+ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__a21o_1
X_15297_ clknet_leaf_17_i_clk _00842_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold307 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14248_ _07050_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold329 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\] VGND VGND VPWR VPWR
+ net446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14179_ _06928_ net293 _06989_ _06990_ _01456_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__o221a_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _01474_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__buf_4
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _01865_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _02195_
+ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07622_ _01303_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
X_07553_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _01249_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07484_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _01122_ _01116_
+ _01047_ _01072_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09223_ _02674_ _02682_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09154_ _02611_ _02615_ _02622_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__or3b_1
XFILLER_0_17_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08105_ _01562_ _01698_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09085_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _02561_
+ _02562_ _02414_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o221a_1
XFILLER_0_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08036_ _01463_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[7\] _01460_ _01634_
+ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09987_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03357_ VGND
+ VGND VPWR VPWR _03358_ sky130_fd_sc_hd__xnor2_1
X_08938_ _02313_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02427_
+ _02428_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08869_ _02329_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _02368_ _02370_ _02309_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__o221a_1
X_10900_ _04153_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nand2_1
X_11880_ _04754_ _05008_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__or3_1
X_10831_ _04077_ _04079_ _04087_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13550_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _06451_ sky130_fd_sc_hd__inv_2
X_10762_ _04023_ net463 _04031_ _04032_ _03814_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12501_ _04538_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13481_ _06210_ net336 _06203_ _06391_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__o211a_1
X_10693_ _03958_ _03956_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__or3_1
X_15220_ clknet_leaf_15_i_clk _00765_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12432_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05489_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15151_ clknet_leaf_125_i_clk _00696_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12363_ _05423_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__buf_2
XFILLER_0_90_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14102_ _06902_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__clkbuf_4
X_11314_ _04503_ _04506_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15082_ clknet_leaf_119_i_clk _00627_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_12294_ _05000_ _05365_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14033_ _06555_ _06867_ _06868_ _06747_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__o211a_1
X_11245_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _04451_ VGND
+ VGND VPWR VPWR _04452_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11176_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__or2_1
X_10127_ _03290_ net503 VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__or2_1
X_14935_ clknet_leaf_110_i_clk net241 VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10058_ _03420_ _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_14_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_14866_ clknet_leaf_84_i_clk _00411_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_13817_ _06663_ _06665_ _06673_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14797_ clknet_leaf_71_i_clk _00342_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_13748_ _06561_ net597 _06485_ _06620_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13679_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _06562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15418_ clknet_leaf_25_i_clk _00963_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15349_ clknet_leaf_29_i_clk _00894_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold104 _00879_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold115 diff3\[5\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold126 net103 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold159 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _03287_ VGND
+ VGND VPWR VPWR _03288_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09841_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _03227_
+ _03229_ _03201_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__a31o_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _03170_ _03171_ _03172_ _03173_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__o31a_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\] _02243_ VGND VGND VPWR
+ VPWR _02244_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\] _02170_ _01879_ VGND
+ VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o21a_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ r_i_alpha1\[7\] _01289_ _01276_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\] _02113_ _02101_ VGND
+ VGND VPWR VPWR _02119_ sky130_fd_sc_hd__a21bo_1
X_07536_ _01240_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07467_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _01081_ _01085_
+ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09206_ _02608_ _02627_ _02651_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07398_ _01076_ _01131_ _01135_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09137_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__or4_4
XFILLER_0_60_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09068_ _02524_ _02543_ _02546_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08019_ _01603_ _01600_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11030_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04270_ VGND
+ VGND VPWR VPWR _04271_ sky130_fd_sc_hd__xnor2_2
X_12981_ _05652_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__and2_1
X_14720_ clknet_leaf_53_i_clk net448 VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11932_ _05020_ _05030_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _04989_ _04987_ _04993_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__o21bai_2
X_14651_ clknet_leaf_49_i_clk _00196_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04075_ VGND
+ VGND VPWR VPWR _04077_ sky130_fd_sc_hd__nand2_1
X_13602_ _06496_ _06497_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__and2b_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _04931_ _04932_ _04786_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__o21ai_1
X_14582_ clknet_leaf_40_i_clk _00127_ VGND VGND VPWR VPWR diff3\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10745_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND VPWR
+ VPWR _04018_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13533_ _06434_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND
+ VGND VPWR VPWR _06436_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13464_ _06374_ _06373_ _06375_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10676_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03943_ VGND
+ VGND VPWR VPWR _03966_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15203_ clknet_leaf_0_i_clk _00748_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12415_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] net653 _05430_ VGND
+ VGND VPWR VPWR _05475_ sky130_fd_sc_hd__o41a_1
X_13395_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06314_ VGND
+ VGND VPWR VPWR _06315_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15134_ clknet_leaf_125_i_clk _00679_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12346_ _05387_ _05398_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15065_ clknet_leaf_102_i_clk _00610_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12277_ _05350_ _05351_ _01250_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14016_ _06851_ _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__xnor2_1
X_11228_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _04420_ _04414_
+ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__a41o_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _04377_ net175 _04219_ _04383_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__o211a_1
X_14918_ clknet_leaf_87_i_clk _00463_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14849_ clknet_leaf_68_i_clk _00394_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[9\] _01916_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[10\]
+ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07321_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ _01048_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__or3_4
XFILLER_0_129_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07252_ net363 net8 _01000_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09824_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _03212_
+ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__or2_1
X_09755_ _03155_ _03157_ _03153_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__a21oi_1
X_08706_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\] _02221_ _02227_ VGND
+ VGND VPWR VPWR _02228_ sky130_fd_sc_hd__o21a_1
X_09686_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _03096_ sky130_fd_sc_hd__or2_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _01864_ _02164_ _02165_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__or3_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _02091_ _02094_ _02086_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07519_ net319 VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08499_ _02014_ _02017_ _02030_ _02040_ _02029_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10530_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _03832_ VGND
+ VGND VPWR VPWR _03833_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10461_ _03772_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12200_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05279_ VGND
+ VGND VPWR VPWR _05285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13180_ _06103_ _06104_ _06097_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__nor3b_1
X_10392_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__or4_1
X_12131_ _05220_ _05221_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12062_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__clkbuf_4
Xhold490 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND VGND VPWR
+ VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ _04254_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12964_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05941_ VGND
+ VGND VPWR VPWR _05942_ sky130_fd_sc_hd__xnor2_1
X_14703_ clknet_leaf_62_i_clk _00248_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11915_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _05041_ _04757_
+ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__mux2_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _05862_ VGND VGND
+ VPWR VPWR _05884_ sky130_fd_sc_hd__and4_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14634_ clknet_leaf_45_i_clk _00179_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _03619_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__clkbuf_4
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04917_ _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__nand2_1
X_14565_ clknet_leaf_35_i_clk _00111_ VGND VGND VPWR VPWR diff2\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10728_ _03995_ net234 _04003_ _04006_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__o211a_1
X_13516_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14496_ clknet_leaf_4_i_clk _00042_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10659_ _03948_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_8_i_clk clknet_4_2_0_i_clk VGND VGND VPWR VPWR clknet_leaf_8_i_clk sky130_fd_sc_hd__clkbuf_16
X_13447_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _06337_ VGND
+ VGND VPWR VPWR _06362_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13378_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _06299_ VGND
+ VGND VPWR VPWR _06300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15117_ clknet_leaf_113_i_clk _00662_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12329_ _05379_ _05398_ _05387_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15048_ clknet_leaf_112_i_clk net144 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_07870_ _01328_ _01487_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__or2_1
X_09540_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ _02918_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__or4_4
X_09471_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02899_ _02900_
+ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08422_ _01962_ _01966_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08353_ _01909_ _01911_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07304_ _01017_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_4
X_08284_ _01330_ _01771_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07235_ _00996_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09807_ _03196_ _03198_ _03199_ _03201_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__a31o_1
X_07999_ net33 net51 VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__and2_1
X_09738_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03142_ VGND
+ VGND VPWR VPWR _03143_ sky130_fd_sc_hd__xnor2_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03079_ VGND
+ VGND VPWR VPWR _03080_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _04848_ _03118_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__and2b_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _05648_ VGND
+ VGND VPWR VPWR _05700_ sky130_fd_sc_hd__xor2_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11631_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _04778_
+ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__nand2_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11562_ _04735_ _04736_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14350_ _07128_ _07130_ _07137_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__nor3_1
XFILLER_0_147_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10513_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _03796_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__o21a_1
X_13301_ _06234_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14281_ _07076_ _07077_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__or2b_1
X_11493_ _04669_ _04673_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13232_ _06178_ _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__nand2_1
X_10444_ _03755_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ _06103_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10375_ _03692_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12114_ _05153_ net424 _05206_ _05207_ _05170_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__o221a_1
X_13094_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _06010_ VGND
+ VGND VPWR VPWR _06057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12045_ _05148_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13996_ _06822_ _06835_ _06829_ _06804_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__or4b_1
XFILLER_0_99_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12947_ _05927_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__buf_2
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _05868_
+ _05845_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ clknet_leaf_44_i_clk _00162_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11829_ _04538_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__clkbuf_4
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14548_ clknet_leaf_40_i_clk _00094_ VGND VGND VPWR VPWR diff1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14479_ clknet_leaf_25_i_clk _00025_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08971_ _02452_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07922_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] _01531_ VGND VGND
+ VPWR VPWR _01532_ sky130_fd_sc_hd__nor2_1
Xhold19 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _01251_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07784_ net232 _01338_ _01420_ _01422_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__o22a_1
X_09523_ _02497_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_109_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_109_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09454_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _02884_ VGND
+ VGND VPWR VPWR _02886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08405_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND VPWR
+ VPWR _01956_ sky130_fd_sc_hd__inv_2
X_09385_ _02308_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08336_ _01893_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR _01898_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08267_ _01750_ _01840_ _01470_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08198_ _01717_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\] _01635_ _01784_
+ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10160_ _03190_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND
+ VGND VPWR VPWR _03514_ sky130_fd_sc_hd__or2_1
X_10091_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _03450_ VGND
+ VGND VPWR VPWR _03451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13850_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _06707_ VGND
+ VGND VPWR VPWR _06708_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12801_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _05789_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__o41a_1
X_10993_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _04237_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13781_ _06643_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__and2b_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _05745_ VGND
+ VGND VPWR VPWR _05746_ sky130_fd_sc_hd__and2_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _05684_ _05685_ _05492_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__and3b_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _07181_ _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11614_ _04774_ _04775_ _04445_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15382_ clknet_leaf_38_i_clk _00927_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12594_ _05615_ _05624_ _04961_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14333_ _01862_ _01032_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__nor2_1
X_11545_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04692_ VGND
+ VGND VPWR VPWR _04722_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11476_ _04659_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__clkbuf_1
X_14264_ _06907_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND
+ VGND VPWR VPWR _07064_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13215_ _06160_ _06163_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__nand2_1
X_10427_ _03724_ _03726_ _03734_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__a31oi_2
X_14195_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _07002_ VGND
+ VGND VPWR VPWR _07003_ sky130_fd_sc_hd__xnor2_2
X_13146_ _06100_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__nor2_2
X_10358_ _03623_ _03677_ _03678_ _03515_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _05652_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__and2_1
X_10289_ net158 _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__or2_1
X_12028_ net169 _05132_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_26_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13979_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06807_ VGND
+ VGND VPWR VPWR _06821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09170_ _02441_ _02629_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08121_ _01691_ _01703_ _01690_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08052_ _01556_ _01642_ _01648_ _01649_ _01485_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08954_ _02342_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__nand2_1
X_07905_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[11\] _01517_ VGND VGND
+ VPWR VPWR _01518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08885_ _01959_ _02383_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__a21bo_1
X_07836_ _01455_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_4
X_07767_ _01412_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
X_09506_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _02932_ VGND
+ VGND VPWR VPWR _02933_ sky130_fd_sc_hd__xor2_2
X_07698_ net340 _01362_ _01358_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _02870_ _01979_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__and2b_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09368_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _02806_
+ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08319_ _01882_ _01883_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__xnor2_1
X_09299_ _02748_ net210 _02749_ _02753_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11330_ _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11261_ _04466_ _03118_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__and2b_1
X_13000_ _05960_ _05974_ _05964_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__a21o_1
X_10212_ _03558_ _03560_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__or2_1
X_11192_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _04394_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__or3_1
X_10143_ _03494_ _03496_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14951_ clknet_leaf_106_i_clk _00496_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10074_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _03410_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13902_ _06501_ _06753_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__and2_1
X_14882_ clknet_leaf_110_i_clk _00427_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13833_ _06563_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _06692_
+ _06693_ _06631_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13764_ _06293_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _06625_ _06633_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__a31o_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10976_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _04221_ VGND
+ VGND VPWR VPWR _04222_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12715_ _05652_ _05730_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13695_ _06565_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _06574_ _06575_ _06526_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__o221a_1
X_15434_ clknet_leaf_27_i_clk _00979_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12646_ _05668_ _05669_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15365_ clknet_leaf_21_i_clk _00910_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12577_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _05607_ VGND
+ VGND VPWR VPWR _05609_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14316_ _07100_ _07108_ _04961_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__o21a_1
X_11528_ _04705_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_10_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15296_ clknet_leaf_14_i_clk net612 VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold308 diff3\[7\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 _00769_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ _07049_ _01512_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__and2b_1
X_11459_ _04640_ _04643_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06985_
+ _06988_ _01862_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__o31ai_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13129_ _06081_ _06075_ _06087_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and3_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08670_ _02194_ _02189_ _02190_ _01868_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__o31a_1
XFILLER_0_89_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07621_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\] _01302_ _01282_
+ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07552_ net413 VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
X_07483_ _01022_ _01114_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__nor2_1
X_09222_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02685_ VGND
+ VGND VPWR VPWR _02686_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09153_ _02611_ _02615_ _02622_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08104_ _01691_ _01697_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09084_ _02552_ _02548_ _02560_ _02369_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08035_ _01465_ _01633_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09986_ _03206_ _03356_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08937_ _02420_ _02421_ _02426_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__o31a_1
X_08868_ _02367_ _02364_ _02366_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__a31o_1
X_07819_ _01447_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
X_08799_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _02312_ sky130_fd_sc_hd__inv_2
X_10830_ _04091_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10761_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _04030_
+ _03997_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__o21ai_1
X_12500_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05541_
+ _05490_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10692_ _03967_ _03972_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__or2_1
X_13480_ _06389_ _06390_ _06232_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12431_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15150_ clknet_leaf_125_i_clk _00695_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ _05234_ _05428_ _05429_ _05343_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14101_ _06923_ _06924_ net358 VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__a21oi_1
X_11313_ _04512_ _04513_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15081_ clknet_leaf_119_i_clk _00626_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_12293_ _05000_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11244_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _04450_ VGND
+ VGND VPWR VPWR _04451_ sky130_fd_sc_hd__xnor2_1
X_14032_ _06562_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _06868_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11175_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
X_10126_ _03476_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__xor2_1
X_14934_ clknet_leaf_108_i_clk _00479_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10057_ _03403_ _03421_ _03412_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14865_ clknet_leaf_84_i_clk _00410_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_13816_ _01765_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14796_ clknet_leaf_71_i_clk _00341_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13747_ _06563_ _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__nand2_1
X_10959_ _04204_ _04207_ _03993_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13678_ _06557_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__clkbuf_4
X_15417_ clknet_leaf_27_i_clk _00962_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12629_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _05640_ VGND
+ VGND VPWR VPWR _05656_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15348_ clknet_leaf_48_i_clk _00893_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold105 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 net110 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ clknet_leaf_51_i_clk _00824_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold127 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold138 net78 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _03227_ _03229_ net395 VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__a21oi_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03151_ VGND
+ VGND VPWR VPWR _03173_ sky130_fd_sc_hd__xor2_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[12\] _02242_ VGND VGND VPWR
+ VPWR _02243_ sky130_fd_sc_hd__xor2_1
X_08653_ _01867_ _02179_ _02180_ _01552_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07604_ diff2\[7\] _01270_ _01272_ diff3\[7\] _01288_ VGND VGND VPWR VPWR _01289_
+ sky130_fd_sc_hd__a221o_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08584_ _01877_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07535_ net381 net346 _01234_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07466_ _01044_ net335 _01192_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09205_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__or2_1
X_07397_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _01080_ _01081_
+ _01134_ _01085_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09136_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _02607_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09067_ _02544_ _02535_ _02545_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08018_ net34 net52 VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09969_ _03341_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__clkbuf_1
X_12980_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05956_ _05844_
+ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__mux2_1
X_11931_ _05029_ _05044_ _05039_ _05052_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__a41oi_2
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ clknet_leaf_50_i_clk net160 VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11862_ _04990_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__xnor2_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06488_ VGND
+ VGND VPWR VPWR _06497_ sky130_fd_sc_hd__nand2_1
X_10813_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04075_ VGND
+ VGND VPWR VPWR _04076_ sky130_fd_sc_hd__or2_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14581_ clknet_leaf_41_i_clk _00126_ VGND VGND VPWR VPWR diff3\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04931_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__and2_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13532_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _06434_ VGND
+ VGND VPWR VPWR _06435_ sky130_fd_sc_hd__and2b_1
X_10744_ _04011_ net562 _04016_ _04017_ _03814_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13463_ _06373_ _06374_ _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10675_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03944_ VGND
+ VGND VPWR VPWR _03965_ sky130_fd_sc_hd__nand2_1
X_15202_ clknet_leaf_0_i_clk _00747_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12414_ _05472_ _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13394_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06235_ VGND VGND
+ VPWR VPWR _06314_ sky130_fd_sc_hd__o31a_1
X_15133_ clknet_leaf_125_i_clk _00678_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12345_ _05140_ net327 _05141_ _05413_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15064_ clknet_leaf_117_i_clk _00609_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12276_ _05344_ _05349_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__and2_1
X_14015_ _06839_ _06842_ _06852_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__a21oi_1
X_11227_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04432_
+ _04414_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__o21a_1
X_11158_ net151 _04379_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ _03035_ _03466_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__nor2_1
X_11089_ _04324_ _03669_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__mux2_1
X_14917_ clknet_leaf_87_i_clk _00462_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14848_ clknet_leaf_85_i_clk _00393_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14779_ clknet_leaf_75_i_clk _00324_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07320_ _01044_ net168 _01065_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07251_ _01005_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09823_ _03184_ net496 _03215_ _03058_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__o211a_1
X_09754_ _03153_ _03155_ _03157_ _02745_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__a31o_1
X_08705_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\] _02221_ _02211_ VGND
+ VGND VPWR VPWR _02227_ sky130_fd_sc_hd__a21bo_1
X_09685_ _03090_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__xnor2_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _02157_ _02150_ _02163_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__a21oi_2
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _02101_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07518_ net67 net318 _01013_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08498_ _02011_ _02028_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07449_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _01159_ _01178_
+ _01179_ _01059_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10460_ _03535_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09119_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out _02591_ VGND
+ VGND VPWR VPWR _02592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10391_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR
+ VPWR _03708_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12130_ _05128_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12061_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _05163_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold480 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold491 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ _04250_ _04253_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__nand2_1
X_12963_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _05941_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14702_ clknet_leaf_62_i_clk _00247_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_11914_ _05038_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__xnor2_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _05871_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _05882_ _05883_ _05751_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__o221a_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ clknet_leaf_58_i_clk _00178_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _04769_ _04977_ _04978_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__a21oi_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ clknet_leaf_40_i_clk _00110_ VGND VGND VPWR VPWR diff2\[8\] sky130_fd_sc_hd__dfxtp_1
X_11776_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _04915_ _04916_
+ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__nand3_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13515_ _06201_ _06419_ _06420_ _06110_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10727_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _03999_
+ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__or2_1
X_14495_ clknet_leaf_5_i_clk _00041_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13446_ _06323_ _06357_ _06358_ _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__a31oi_2
X_10658_ _03925_ _03927_ _03937_ _03949_ _03936_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__o32a_1
XFILLER_0_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13377_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06298_ VGND
+ VGND VPWR VPWR _06299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10589_ _03605_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _03885_
+ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15116_ clknet_leaf_113_i_clk _00661_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12328_ _05383_ _05385_ _05382_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15047_ clknet_leaf_102_i_clk _00592_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
X_12259_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05336_ _01249_
+ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__mux2_1
X_09470_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02899_ _02885_
+ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__a21o_1
X_08421_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\] _01965_ VGND VGND VPWR
+ VPWR _01969_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08352_ _01909_ _01911_ _01866_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07303_ _01047_ _01048_ _01049_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08283_ _01454_ _01849_ _01854_ _01855_ _01766_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__o311a_1
XFILLER_0_116_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07234_ net353 net17 _00993_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09806_ _03182_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07998_ _01597_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__and2_1
X_09737_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03141_ VGND
+ VGND VPWR VPWR _03142_ sky130_fd_sc_hd__xor2_2
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09668_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _03069_ _02770_
+ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__o21a_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _02146_ _02148_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__xnor2_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _02754_ net478 _02749_ _03016_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__o211a_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _04775_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__or3_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11561_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04723_ _04732_
+ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13300_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _06234_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10512_ _03792_ _03797_ _03807_ _03811_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14280_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _07023_ VGND
+ VGND VPWR VPWR _07077_ sky130_fd_sc_hd__or2_1
X_11492_ _04669_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13231_ _06177_ _06172_ _06174_ _05844_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10443_ _03743_ _03749_ _03747_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ _06104_ _06107_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10374_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _03691_ VGND
+ VGND VPWR VPWR _03693_ sky130_fd_sc_hd__nor2_1
X_12113_ _05205_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _05129_
+ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__a21o_1
X_13093_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06010_ _06053_
+ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__a21o_1
X_12044_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND VPWR
+ VPWR _05149_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13995_ _06811_ _06816_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12946_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _05927_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12877_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _05868_
+ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__and2_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ clknet_leaf_42_i_clk _00161_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_11828_ _04956_ _04958_ _04962_ _04758_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__o31ai_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14547_ clknet_leaf_41_i_clk _00093_ VGND VGND VPWR VPWR diff1\[6\] sky130_fd_sc_hd__dfxtp_1
X_11759_ _04853_ _04856_ _04888_ _04881_ _04897_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14478_ clknet_leaf_7_i_clk _00024_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13429_ _06338_ _06344_ _06345_ _06199_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08970_ _02448_ _02453_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__and2_1
X_07921_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[13\]
+ _01522_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__and3_1
X_07852_ _01472_ _01468_ _01469_ _01453_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__a31o_1
Xinput1 i_rst_n VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_07783_ _01338_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09522_ _02746_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02946_
+ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09453_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _02884_ VGND
+ VGND VPWR VPWR _02885_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08404_ _01891_ net531 _01954_ _01955_ _01908_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09384_ _02824_ _02822_ _02823_ _02761_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08335_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[5\] _01892_ VGND VGND
+ VPWR VPWR _01897_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08266_ _01750_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08197_ _01330_ _01568_ _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10090_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _03449_ VGND
+ VGND VPWR VPWR _03450_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_7_i_clk sky130_fd_sc_hd__clkbuf_16
X_12800_ _05783_ _05788_ _05795_ _05801_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__and4_1
X_13780_ _06646_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__clkbuf_4
X_10992_ _04236_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _05744_ VGND
+ VGND VPWR VPWR _05745_ sky130_fd_sc_hd__xor2_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12662_ _05683_ _05680_ _05682_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__or3_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _07156_ VGND
+ VGND VPWR VPWR _07182_ sky130_fd_sc_hd__nand2_1
X_11613_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__or2_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15381_ clknet_leaf_38_i_clk _00926_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12593_ _05622_ _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14332_ _06910_ net423 _01766_ _07121_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__o211a_1
X_11544_ _04390_ net504 _04387_ _04721_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14263_ _07061_ _07062_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11475_ _04468_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13214_ _06160_ _06163_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10426_ _03738_ _03733_ _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14194_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _07001_ VGND
+ VGND VPWR VPWR _07002_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13145_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06101_ VGND
+ VGND VPWR VPWR _06102_ sky130_fd_sc_hd__xnor2_1
X_10357_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _03678_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06041_ _05844_
+ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__mux2_1
X_10288_ _03608_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__buf_2
X_12027_ _05130_ net162 _04979_ _05136_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__o211a_1
X_13978_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06807_ VGND
+ VGND VPWR VPWR _06820_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12929_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05912_
+ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08120_ _01562_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08051_ _01625_ _01638_ _01646_ _01572_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__or4_4
X_07904_ _01515_ _01516_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\]
+ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__mux2_1
X_08884_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _02371_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07835_ _01454_ net242 _01456_ _01459_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07766_ net438 _01410_ _01411_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__mux2_1
X_09505_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02918_ _02771_
+ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07697_ _01360_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _02746_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02868_
+ _02869_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__a22oi_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09367_ _02757_ net580 _02810_ _02811_ _02689_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08318_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\]
+ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__xor2_2
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09298_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _02751_
+ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08249_ _01465_ _01826_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11260_ _04396_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04464_
+ _04465_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_104_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10211_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03559_ VGND
+ VGND VPWR VPWR _03560_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11191_ _04390_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _04405_ _04406_ _04360_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10142_ _03494_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nor2_1
X_14950_ clknet_leaf_107_i_clk _00495_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10073_ _03412_ _03421_ _03434_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__or3b_1
X_13901_ _06751_ _06752_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _06554_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__a2bb2o_1
X_14881_ clknet_leaf_110_i_clk net131 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13832_ _06685_ _06688_ _06691_ _06584_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_97_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13763_ _06293_ _06632_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__nor2_1
X_10975_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _04220_ VGND
+ VGND VPWR VPWR _04221_ sky130_fd_sc_hd__xnor2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _05729_ _05489_
+ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13694_ _06568_ _06573_ _06555_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__a21o_1
X_15433_ clknet_leaf_28_i_clk _00978_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_12645_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _05648_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__o41a_2
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15364_ clknet_leaf_23_i_clk _00909_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12576_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _05607_ VGND
+ VGND VPWR VPWR _05608_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14315_ _07106_ _07107_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11527_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04692_ VGND
+ VGND VPWR VPWR _04706_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15295_ clknet_leaf_19_i_clk _00840_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14246_ _06903_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _07047_
+ _07048_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__a22oi_1
Xhold309 diff3\[14\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ _04631_ _04635_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10409_ _03705_ _03714_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14177_ _06985_ _06988_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__o21a_1
X_11389_ _04581_ _04577_ _04578_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_108_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_108_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _06085_ _06086_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__or2_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _06005_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07620_ r_i_alpha1\[10\] _01301_ _01276_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07551_ net66 net412 _01012_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07482_ _01095_ net369 _01203_ _01204_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09221_ _02544_ _02684_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09152_ _02620_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08103_ _01641_ _01692_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09083_ _02552_ _02548_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08034_ _01630_ _01632_ _01470_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09985_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _03315_ _03355_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__or4_4
XFILLER_0_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08936_ _02420_ _02421_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_72_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08867_ _02313_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__buf_4
X_07818_ net396 _01446_ _00992_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__mux2_1
X_08798_ _02311_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_87_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07749_ _01398_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10760_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _04030_
+ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09419_ _02595_ net449 _02747_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_i_clk clknet_4_2_0_i_clk VGND VGND VPWR VPWR clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10691_ _03977_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12430_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12361_ _05139_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _05429_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14100_ _06646_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ _06914_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__or3_1
X_11312_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _04511_ VGND
+ VGND VPWR VPWR _04513_ sky130_fd_sc_hd__and2b_1
X_15080_ clknet_leaf_120_i_clk _00625_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_25_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12292_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05364_ VGND
+ VGND VPWR VPWR _05365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14031_ _06863_ _06866_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11243_ _04061_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND
+ VGND VPWR VPWR _04450_ sky130_fd_sc_hd__and2b_1
X_11174_ _04390_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _04387_ _04392_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__o211a_1
X_10125_ _03480_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nand2_1
X_14933_ clknet_leaf_106_i_clk _00478_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
X_10056_ _03394_ _03413_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__nor2_1
X_14864_ clknet_leaf_85_i_clk _00409_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13815_ _06677_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
X_14795_ clknet_leaf_68_i_clk _00340_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13746_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _06618_
+ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__xnor2_1
X_10958_ _04177_ _04205_ _04206_ _04179_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13677_ _06556_ net288 _06485_ _06560_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10889_ _04142_ _04144_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12628_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _05641_ VGND
+ VGND VPWR VPWR _05655_ sky130_fd_sc_hd__nand2_1
X_15416_ clknet_leaf_27_i_clk _00961_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15347_ clknet_leaf_38_i_clk _00892_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12559_ _05579_ _05583_ _05580_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold106 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
X_15278_ clknet_leaf_51_i_clk net296 VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold117 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _06907_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND
+ VGND VPWR VPWR _07034_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_8_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_09770_ _03155_ _03169_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\] _02231_ _01880_ VGND
+ VGND VPWR VPWR _02242_ sky130_fd_sc_hd__o21a_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _01873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _02180_ sky130_fd_sc_hd__or2_1
X_07603_ _01273_ diff1\[7\] VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08583_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] VGND VGND VPWR
+ VPWR _02117_ sky130_fd_sc_hd__inv_2
X_07534_ _01239_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07465_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _01159_ _01190_
+ _01191_ _01030_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09204_ _02333_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND
+ VGND VPWR VPWR _02669_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07396_ _01132_ _01133_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09135_ _02606_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09066_ _02544_ _02535_ _02528_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08017_ _01613_ _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__xnor2_1
X_09968_ _03024_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__and2_1
X_08919_ _02152_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _02412_ sky130_fd_sc_hd__nor2_1
X_09899_ _03237_ net526 _03278_ _03279_ _03258_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__o221a_1
X_11930_ _05036_ _05049_ _05050_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__a21oi_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04991_ VGND
+ VGND VPWR VPWR _04992_ sky130_fd_sc_hd__xnor2_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06488_ VGND
+ VGND VPWR VPWR _06496_ sky130_fd_sc_hd__nor2_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10812_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _04074_ VGND
+ VGND VPWR VPWR _04075_ sky130_fd_sc_hd__xnor2_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ clknet_leaf_39_i_clk _00125_ VGND VGND VPWR VPWR diff3\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _04925_ _04927_ _04923_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06433_ VGND
+ VGND VPWR VPWR _06434_ sky130_fd_sc_hd__xnor2_1
X_10743_ _03669_ _04014_ _04015_ _03994_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13462_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _06351_ VGND
+ VGND VPWR VPWR _06375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10674_ _03625_ net408 _03620_ _03964_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15201_ clknet_leaf_1_i_clk _00746_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12413_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05430_ VGND
+ VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13393_ _06313_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15132_ clknet_leaf_122_i_clk _00677_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12344_ _05142_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15063_ clknet_leaf_117_i_clk _00608_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12275_ _05344_ _05349_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__nor2_1
X_14014_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _06845_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__o21a_1
X_11226_ _04431_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _04435_ _04436_ _04360_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11157_ _04377_ net223 _04219_ _04382_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__o211a_1
X_10108_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _03465_ VGND
+ VGND VPWR VPWR _03466_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11088_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04313_ _04034_
+ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__o21a_1
X_14916_ clknet_leaf_87_i_clk _00461_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10039_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _03406_ sky130_fd_sc_hd__or2_1
X_14847_ clknet_leaf_86_i_clk _00392_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14778_ clknet_leaf_76_i_clk _00323_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13729_ _06561_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _06485_ _06604_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07250_ net354 net7 _01000_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09822_ net254 _03190_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09753_ _03138_ _03156_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__nand2_1
X_08704_ _02022_ net581 _02225_ _02226_ _02055_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__o221a_1
X_09684_ _03054_ _03063_ _03074_ _03083_ _03093_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__a41o_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _02157_ _02150_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__and3_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\] _02100_ VGND VGND VPWR
+ VPWR _02102_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07517_ _01230_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08497_ _02037_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07448_ _01010_ _01020_ _01022_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07379_ _01044_ net182 _01118_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09118_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _02591_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10390_ _03623_ _03706_ _03707_ _03515_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09049_ _02528_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12060_ _05153_ net525 _05161_ _05162_ _04965_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__o221a_1
Xhold470 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND VGND VPWR
+ VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _04250_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__or2_1
Xhold492 net87 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
X_12962_ _05931_ _05935_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11913_ _05021_ _05039_ _05029_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__o21a_1
X_14701_ clknet_leaf_62_i_clk _00246_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12893_ _05881_ _05879_ _05880_ _05860_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__a31o_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _04786_ net414 _01794_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__o21ai_1
X_14632_ clknet_leaf_58_i_clk _00177_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ clknet_leaf_40_i_clk _00109_ VGND VGND VPWR VPWR diff2\[7\] sky130_fd_sc_hd__dfxtp_1
X_11775_ _04915_ _04916_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10726_ _03995_ net265 _04003_ _04005_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__o211a_1
X_13514_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _06420_ sky130_fd_sc_hd__or2_1
X_14494_ clknet_leaf_4_i_clk _00040_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13445_ _06339_ _06359_ _06358_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10657_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03934_ _03923_
+ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10588_ _03872_ _03878_ _03884_ _03605_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12327_ _05395_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__or2_1
X_15115_ clknet_leaf_112_i_clk _00660_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15046_ clknet_leaf_98_i_clk _00591_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12258_ _05332_ _05335_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11209_ _04421_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__inv_2
X_12189_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR _05275_ sky130_fd_sc_hd__inv_2
X_08420_ _01867_ _01967_ _01968_ _01552_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08351_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[7\] _01903_ _01910_
+ _01550_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__a22o_1
X_07302_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _01033_ VGND
+ VGND VPWR VPWR _01049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08282_ _01464_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[16\] VGND VGND VPWR
+ VPWR _01855_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07233_ _00995_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09805_ _03198_ _03199_ _03196_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__a21oi_1
X_07997_ net52 net34 VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__or2b_2
X_09736_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03130_ _02772_
+ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09667_ _03078_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\] _02147_ VGND VGND VPWR
+ VPWR _02148_ sky130_fd_sc_hd__xnor2_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _03014_ _03015_ _02755_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__o21ai_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[12\] _02085_ VGND VGND VPWR
+ VPWR _02087_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11560_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04723_ VGND
+ VGND VPWR VPWR _04735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10511_ _03815_ _03816_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11491_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04672_ VGND
+ VGND VPWR VPWR _04673_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13230_ _06172_ _06174_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10442_ _03752_ _03754_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13161_ _06115_ _06116_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__nor2_2
XFILLER_0_60_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10373_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _03691_ VGND
+ VGND VPWR VPWR _03692_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12112_ _05205_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _05206_ sky130_fd_sc_hd__nor2_1
X_13092_ _06049_ _06055_ _04961_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12043_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND VPWR
+ VPWR _05148_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13994_ _06822_ _06833_ _06829_ _06828_ _06821_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__o311a_1
XFILLER_0_99_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12945_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05922_
+ _05921_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__a21oi_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _05567_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _05858_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__o31a_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ clknet_leaf_45_i_clk _00160_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_11827_ _04956_ _04958_ _04962_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__o21a_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _04888_ _04883_ _04897_ _04900_ _04896_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a32o_1
X_14546_ clknet_leaf_41_i_clk _00092_ VGND VGND VPWR VPWR diff1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10709_ _03993_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11689_ _04756_ _04837_ _04838_ _04739_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__o211a_1
X_14477_ clknet_leaf_7_i_clk _00023_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13428_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _06337_ VGND
+ VGND VPWR VPWR _06345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13359_ _04538_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07920_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\] _01528_
+ _01530_ _01513_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__o221a_1
X_15029_ clknet_leaf_103_i_clk _00574_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07851_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] VGND VGND VPWR VPWR
+ _01472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 i_valid_in VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
X_07782_ net15 net14 net16 VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__a21o_1
X_09521_ _02939_ _02945_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _02883_ VGND
+ VGND VPWR VPWR _02884_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08403_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[16\] _01952_ _01953_
+ _01870_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__o31ai_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09383_ _02822_ _02823_ _02824_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08334_ _01891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _01895_ _01896_ _01661_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08265_ _01728_ _01830_ _01839_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08196_ _01470_ _01781_ _01782_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in
+ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09719_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _03125_ VGND
+ VGND VPWR VPWR _03126_ sky130_fd_sc_hd__nand2_1
X_10991_ _03976_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05734_ _05525_
+ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__o21a_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _05680_ _05682_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__o21a_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14400_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _07144_ VGND
+ VGND VPWR VPWR _07181_ sky130_fd_sc_hd__or2_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _05608_ _05616_ _05621_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__a21o_1
X_15380_ clknet_leaf_29_i_clk _00925_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11543_ _04719_ _04720_ _04391_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14331_ _07119_ _07120_ _06904_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14262_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _07042_ _07057_
+ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__a21bo_1
X_11474_ _04656_ _04657_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ _04375_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_150_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13213_ _06161_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__or2_1
X_10425_ _03738_ _03733_ _03722_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__o21ba_1
X_14193_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13144_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06094_ _05878_
+ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__o21a_1
X_10356_ _03672_ _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__xor2_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _06037_ _06040_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__xor2_1
X_10287_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__clkbuf_4
X_12026_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] _05132_
+ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ _06555_ _06818_ _06819_ _06747_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12928_ _05567_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05904_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__o31a_1
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__clkbuf_4
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14529_ clknet_leaf_39_i_clk _00075_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08050_ _01638_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08952_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _02441_ sky130_fd_sc_hd__inv_2
X_07903_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\] _01508_ VGND VGND
+ VPWR VPWR _01516_ sky130_fd_sc_hd__nand2_1
X_08883_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _02376_
+ _01958_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__a21oi_1
X_07834_ net159 _01457_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__or2_1
X_07765_ _00992_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__buf_4
X_09504_ _02754_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02749_
+ _02931_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07696_ net5 _01003_ _01355_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__or3_2
XFILLER_0_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09435_ _02861_ _02862_ _02867_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o31a_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09366_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _02809_
+ _02755_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08317_ _01881_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__buf_4
X_09297_ _02748_ net174 _02749_ _02752_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08248_ _01684_ _01825_ _01329_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08179_ net28 net46 VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nand2_1
X_10210_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _03536_ _03207_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__o31a_1
X_11190_ net622 _04404_ _04391_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__o21ai_1
X_10141_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03495_ VGND
+ VGND VPWR VPWR _03496_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10072_ _03414_ _03434_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__nand2_1
X_13900_ _06749_ _06750_ _06748_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__o21a_1
X_14880_ clknet_leaf_110_i_clk net137 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13831_ _06685_ _06688_ _06691_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10974_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13762_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06627_
+ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _05726_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13693_ _06568_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15432_ clknet_leaf_28_i_clk _00977_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_12644_ _05643_ _05647_ _05657_ _05663_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12575_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05606_ VGND
+ VGND VPWR VPWR _05607_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15363_ clknet_leaf_21_i_clk _00908_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14314_ _07080_ _07105_ _07102_ _07104_ _06926_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__a41o_1
X_11526_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04692_ VGND
+ VGND VPWR VPWR _04705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15294_ clknet_leaf_17_i_clk net468 VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11457_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _04641_ VGND
+ VGND VPWR VPWR _04642_ sky130_fd_sc_hd__nand2_1
X_14245_ _07046_ _07040_ _07043_ _01861_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__o31a_1
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10408_ _03722_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14176_ _06647_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__xor2_1
X_11388_ _04577_ _04578_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _06082_ _06084_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__and2_1
X_10339_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _03658_
+ _03651_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__o21a_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _06009_ _06017_ _06021_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__nor3_1
X_12009_ _05116_ _05120_ _05124_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07550_ net433 VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
X_07481_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _01045_ _01088_
+ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09220_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _02671_ _02343_
+ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_4_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09151_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _02619_ VGND
+ VGND VPWR VPWR _02621_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08102_ net23 net41 _01695_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09082_ _02558_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08033_ _01627_ _01631_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09984_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08935_ _02424_ _02425_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08866_ _02364_ _02366_ _02367_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__a21oi_1
X_07817_ net9 _01445_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__xnor2_1
X_08797_ _01870_ _02310_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__and2_1
X_07748_ net394 _01397_ _01358_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07679_ net190 _01345_ _01346_ _01348_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09418_ _02595_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _02854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10690_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03944_ VGND
+ VGND VPWR VPWR _03978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09349_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02790_
+ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12360_ _05426_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11311_ _04511_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _04512_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12291_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05164_ VGND VGND VPWR
+ VPWR _05364_ sky130_fd_sc_hd__o31a_1
X_14030_ _06839_ _06864_ _06865_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__a21oi_2
X_11242_ _04431_ net540 _04448_ _04449_ _04360_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11173_ _04391_ net285 VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10124_ _03283_ _03479_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14932_ clknet_leaf_81_i_clk _00477_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10055_ _03418_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__and2_1
X_14863_ clknet_leaf_85_i_clk _00408_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_13814_ _06501_ _06676_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14794_ clknet_leaf_66_i_clk _00339_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_13745_ _06615_ _06617_ _06587_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__mux2_1
X_10957_ _04184_ _04191_ _04198_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13676_ _06557_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__or2_1
X_10888_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04143_ VGND
+ VGND VPWR VPWR _04144_ sky130_fd_sc_hd__xor2_4
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15415_ clknet_leaf_26_i_clk _00960_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12627_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05648_ _05643_
+ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15346_ clknet_leaf_38_i_clk _00891_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12558_ _05590_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11509_ _04431_ net564 _04688_ _04689_ _04539_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__o221a_1
X_15277_ clknet_leaf_17_i_clk _00822_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12489_ _05500_ net584 _05495_ _05533_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold107 diff2\[6\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _00485_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _00937_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ _07029_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _06972_ _06973_ _06934_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__mux2_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _02047_ _02233_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _02177_ _02178_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__and2b_1
X_07602_ _01287_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
X_08582_ _02022_ net499 _02115_ _02116_ _02055_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07533_ net384 net334 _01234_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__mux2_1
X_07464_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _01122_ _01071_
+ _01047_ _01057_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09203_ _02322_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _02667_
+ _02668_ _02414_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07395_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _01123_ VGND
+ VGND VPWR VPWR _01133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09134_ _02605_ _01979_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09065_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR
+ VPWR _02544_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08016_ _01614_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09967_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03339_ _03185_
+ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__mux2_1
X_08918_ _02321_ _02409_ _02381_ _02411_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__o211a_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _03276_
+ _03277_ _03186_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__o31ai_1
X_08849_ _02321_ net355 _01945_ _02353_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__o211a_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _04794_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__o21a_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _04074_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_95_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11791_ _04557_ _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__xor2_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_107_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_107_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13530_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _06398_
+ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__nor2_1
X_10742_ _04014_ _04015_ _03669_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10673_ _03956_ _03959_ _03631_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a211o_1
X_13461_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _06351_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__o21a_1
X_15200_ clknet_leaf_2_i_clk _00745_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12412_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05430_ VGND
+ VGND VPWR VPWR _05472_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13392_ _06069_ _06312_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__and2_1
X_15131_ clknet_leaf_121_i_clk _00676_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12343_ _05409_ _05411_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15062_ clknet_leaf_117_i_clk _00607_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12274_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _05348_ VGND
+ VGND VPWR VPWR _05349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11225_ net387 _04434_ _04376_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a21o_1
X_14013_ _06849_ _06850_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__and2_1
X_11156_ net122 _04379_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10107_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _03206_ VGND VGND VPWR
+ VPWR _03465_ sky130_fd_sc_hd__o31a_1
X_11087_ _04323_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
X_14915_ clknet_leaf_81_i_clk _00460_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10038_ _03403_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__and2_1
X_14846_ clknet_leaf_85_i_clk _00391_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_14777_ clknet_leaf_76_i_clk _00322_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11989_ _05104_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13728_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06602_
+ _06603_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13659_ _06501_ _06547_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_71_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15329_ clknet_leaf_17_i_clk _00874_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09821_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _03213_
+ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__xnor2_1
X_09752_ _03133_ _03143_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__nor2_1
X_08703_ _02222_ _02224_ _01866_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__a21o_1
X_09683_ _03074_ _03091_ _03083_ _03092_ _03082_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__a32o_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _02161_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\] _02100_ VGND VGND VPWR
+ VPWR _02101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07516_ net371 net245 _01013_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08496_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[8\] _02036_ VGND VGND VPWR
+ VPWR _02038_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07447_ _01010_ _01024_ _01052_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07378_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _01045_ _01115_
+ _01117_ _01059_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09117_ _02585_ _02583_ _02588_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__or3b_1
X_09048_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _02527_ VGND
+ VGND VPWR VPWR _02529_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold460 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04252_ VGND
+ VGND VPWR VPWR _04253_ sky130_fd_sc_hd__xor2_1
Xhold482 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold493 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
X_12961_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _05934_ VGND
+ VGND VPWR VPWR _05939_ sky130_fd_sc_hd__and2_1
X_14700_ clknet_leaf_63_i_clk _00245_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_11912_ _05014_ _05017_ _05028_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__o21ai_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _05879_ _05880_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__a21oi_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ clknet_leaf_42_i_clk _00176_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_11843_ _04975_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__xnor2_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ clknet_leaf_41_i_clk _00108_ VGND VGND VPWR VPWR diff2\[6\] sky130_fd_sc_hd__dfxtp_1
X_11774_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04904_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__or3b_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13513_ _06417_ _06418_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__xnor2_1
X_10725_ net261 _03999_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__or2_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ clknet_leaf_4_i_clk _00039_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13444_ _06327_ _06338_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10656_ _03899_ _03902_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10587_ _03872_ _03878_ _03884_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__a21o_1
X_13375_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _06296_
+ net611 _06285_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__o221a_1
XFILLER_0_106_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15114_ clknet_leaf_112_i_clk _00659_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12326_ _05392_ _05394_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15045_ clknet_leaf_98_i_clk _00590_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12257_ _05309_ _05321_ _05333_ _05334_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11208_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _04407_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__or3_1
X_12188_ _05255_ _05273_ _05265_ _05235_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__or4b_4
X_11139_ _04369_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14829_ clknet_leaf_77_i_clk _00374_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08350_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] _01897_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[7\]
+ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07301_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__or4_4
X_08281_ _01852_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07232_ net332 net16 _00993_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] _03193_
+ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nand2_1
X_07996_ net34 net52 VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__or2b_1
X_09735_ _02748_ _03139_ _03140_ _03058_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__o211a_1
X_09666_ _03024_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\]
+ _01879_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__o21a_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08548_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[12\] _02085_ VGND VGND VPWR
+ VPWR _02086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08479_ _01869_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10510_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03796_ VGND
+ VGND VPWR VPWR _03816_ sky130_fd_sc_hd__nand2_1
X_11490_ _04413_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10441_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03753_ VGND
+ VGND VPWR VPWR _03754_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13160_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06114_ VGND
+ VGND VPWR VPWR _06116_ sky130_fd_sc_hd__nor2_1
X_10372_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03690_ VGND
+ VGND VPWR VPWR _03691_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12111_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND VGND VPWR
+ VPWR _05205_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13091_ _06053_ _06054_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12042_ _05140_ net507 _05146_ _05147_ _04965_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__o221a_1
Xhold290 net62 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13993_ _06809_ _06814_ _06815_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12944_ _05871_ net467 _05924_ _05925_ _05910_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _05566_ _05862_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nand2_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ clknet_leaf_42_i_clk _00159_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_11826_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04930_ VGND
+ VGND VPWR VPWR _04962_ sky130_fd_sc_hd__xnor2_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14545_ clknet_leaf_39_i_clk _00091_ VGND VGND VPWR VPWR diff1\[4\] sky130_fd_sc_hd__dfxtp_1
X_11757_ _04886_ _04895_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__nand2_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _03993_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14476_ clknet_leaf_7_i_clk _00022_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
X_11688_ _04765_ net633 VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13427_ _06339_ _06341_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nand2_1
X_10639_ _03932_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13358_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06282_
+ _06232_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12309_ _05379_ _05380_ _05234_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a21o_1
X_13289_ _05927_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _06214_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15028_ clknet_leaf_96_i_clk _00573_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07850_ _01468_ _01469_ _01470_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__a21oi_1
X_07781_ _00991_ _01334_ net16 VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 in_alpha[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ _02939_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__nand2_1
X_09451_ _02770_ _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__nand2_1
X_08402_ _01952_ _01953_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09382_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR _02824_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08333_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[5\] _01894_ _01877_
+ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08264_ _01838_ _01706_ _01729_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08195_ _01565_ _01780_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07979_ _01579_ _01581_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__xnor2_1
X_09718_ _03109_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__inv_2
X_10990_ _03996_ _04231_ _04232_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09649_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03060_ VGND
+ VGND VPWR VPWR _03062_ sky130_fd_sc_hd__nor2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12660_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05641_ VGND
+ VGND VPWR VPWR _05683_ sky130_fd_sc_hd__xor2_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ _04770_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__clkbuf_4
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12591_ _05608_ _05616_ _05621_ _05486_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14330_ _07113_ _07118_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11542_ _04712_ _04718_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14261_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _07023_ VGND
+ VGND VPWR VPWR _07061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11473_ _04653_ _04655_ _04651_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13212_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _06142_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__o41a_1
X_10424_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR _03738_ sky130_fd_sc_hd__inv_2
X_14192_ _06928_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _06999_
+ _07000_ _01456_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13143_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR _06100_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10355_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _03675_ VGND
+ VGND VPWR VPWR _03676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _06029_ _06038_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__o21a_1
X_10286_ _01251_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__clkbuf_4
X_12025_ _05130_ net209 _04979_ _05135_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13976_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND
+ VGND VPWR VPWR _06819_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12927_ _05566_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05905_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__nand3_1
XFILLER_0_69_860 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12858_ _05844_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__buf_2
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11809_ _04941_ _04944_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12789_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05797_ _05489_
+ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__mux2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14528_ clknet_leaf_42_i_clk _00074_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14459_ clknet_leaf_40_i_clk _00005_ VGND VGND VPWR VPWR r_i_alpha1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08951_ _02424_ _02427_ _02435_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__a21boi_1
Xclkbuf_4_0_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_07902_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\] _01514_ VGND VGND
+ VPWR VPWR _01515_ sky130_fd_sc_hd__or2_1
X_08882_ _01455_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07833_ _01454_ net206 _01456_ _01458_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__o211a_1
X_07764_ _01408_ _01409_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09503_ _02929_ _02930_ _02747_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07695_ net5 _01355_ _01003_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09434_ _02861_ _02862_ _02867_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__o21ai_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09365_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _02809_
+ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08316_ _01880_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__buf_2
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09296_ net145 _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08247_ _01681_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08178_ _01764_ _01767_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10140_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _03477_ _03205_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__o31a_1
XFILLER_0_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10071_ _03420_ _03426_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__and2_1
X_13830_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _06684_ VGND
+ VGND VPWR VPWR _06691_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _06565_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _06629_ _06630_ _06631_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__o221a_1
X_10973_ _03619_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__buf_4
X_12712_ _05727_ _05717_ _05714_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a21o_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _06571_ _06572_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15431_ clknet_leaf_28_i_clk _00976_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_12643_ _05666_ _05667_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15362_ clknet_leaf_21_i_clk _00907_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_12574_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05598_ _05526_
+ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14313_ _07080_ _07102_ _07104_ _07105_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11525_ _04704_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15293_ clknet_leaf_17_i_clk _00838_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14244_ _07040_ _07043_ _07046_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11456_ _04634_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03721_ VGND
+ VGND VPWR VPWR _03723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14175_ _06928_ net278 _06986_ _06987_ _06922_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__o221a_1
X_11387_ _04579_ _04580_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ _06082_ _06084_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__nor2_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _03625_ net428 _03620_ _03662_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__o211a_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06003_ VGND
+ VGND VPWR VPWR _06025_ sky130_fd_sc_hd__xnor2_1
X_10269_ _03607_ net216 _03568_ _03610_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__o211a_1
X_12008_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05081_ VGND
+ VGND VPWR VPWR _05124_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13959_ _06803_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07480_ _01076_ _01110_ _01107_ _01080_ _01202_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09150_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _02619_ VGND
+ VGND VPWR VPWR _02620_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08101_ _01682_ _01694_ _01681_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__a21oi_1
X_09081_ _02555_ _02556_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08032_ _01613_ _01616_ _01610_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput50 in_y[3] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _03352_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08934_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02423_ VGND
+ VGND VPWR VPWR _02425_ sky130_fd_sc_hd__or2_1
X_08865_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR _02367_ sky130_fd_sc_hd__inv_2
X_07816_ net8 _01441_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__or2b_1
X_08796_ _01252_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__buf_4
X_07747_ _01003_ _01395_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07678_ _01344_ _01347_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__nor2_1
X_09417_ _02754_ _02851_ _02749_ _02853_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09279_ _02313_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _02736_
+ _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_7_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11310_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04510_ VGND
+ VGND VPWR VPWR _04511_ sky130_fd_sc_hd__xor2_1
X_12290_ _04996_ _05355_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11241_ _04447_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _04376_
+ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11172_ _04378_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__buf_4
XFILLER_0_101_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10123_ _03283_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__or2_1
X_14931_ clknet_leaf_81_i_clk _00476_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10054_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03410_ VGND
+ VGND VPWR VPWR _03419_ sky130_fd_sc_hd__or2_1
X_14862_ clknet_leaf_85_i_clk _00407_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13813_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _06675_ _06562_
+ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__mux2_1
X_14793_ clknet_leaf_66_i_clk _00338_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13744_ _06616_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__inv_2
X_10956_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13675_ _06556_ net220 _06485_ _06559_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__o211a_1
X_10887_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04108_ _04132_
+ _04035_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__o31a_2
XFILLER_0_128_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15414_ clknet_leaf_26_i_clk _00959_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_12626_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _05648_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15345_ clknet_leaf_48_i_clk _00890_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12557_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05589_ VGND
+ VGND VPWR VPWR _05591_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11508_ _04685_ _04687_ _04376_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15276_ clknet_leaf_17_i_clk _00821_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12488_ _05501_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__nand2_1
Xhold108 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14227_ _07030_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__nand2_1
Xhold119 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11439_ _04623_ _04625_ _04375_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14158_ _06966_ _06968_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__nand2_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _01252_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__clkbuf_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _06913_ _06914_ _06647_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08650_ _02161_ _02165_ _02176_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__or3_1
X_07601_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] _01286_ _01282_ VGND
+ VGND VPWR VPWR _01287_ sky130_fd_sc_hd__mux2_1
X_08581_ _02101_ _02107_ _02114_ _01924_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07532_ net349 VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07463_ _01080_ _01066_ _01067_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09202_ _02664_ _02666_ _02333_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07394_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _01123_ VGND
+ VGND VPWR VPWR _01132_ sky130_fd_sc_hd__or2_4
XFILLER_0_60_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09133_ _02319_ _02595_ _02604_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09064_ _02530_ _02536_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08015_ _01589_ _01593_ _01597_ _01588_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09966_ _03335_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__xnor2_1
X_08917_ _02404_ _02410_ _02314_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a21o_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _03276_ _03277_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__o21a_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08848_ _02322_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__nand2_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _02270_ _02291_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__and2b_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _04065_ _04069_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__nor2_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _04915_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__clkbuf_4
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10741_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13460_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _06352_ _06365_
+ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__o21a_1
X_10672_ _03960_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12411_ _05142_ net565 _05470_ _05471_ _05391_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__o221a_1
X_13391_ _06310_ _06311_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ _06200_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_106_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15130_ clknet_leaf_122_i_clk _00675_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12342_ _05410_ _05399_ _05395_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15061_ clknet_leaf_102_i_clk _00606_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12273_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _05347_ VGND
+ VGND VPWR VPWR _05348_ sky130_fd_sc_hd__xnor2_1
X_14012_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06837_ VGND
+ VGND VPWR VPWR _06850_ sky130_fd_sc_hd__nand2_1
X_11224_ net387 _04434_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__nor2_1
X_11155_ _04377_ net251 _04219_ _04381_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10106_ _03464_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
X_11086_ _03976_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__and2_1
X_14914_ clknet_leaf_81_i_clk _00459_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10037_ _03396_ _03402_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__nand2_1
X_14845_ clknet_leaf_85_i_clk _00390_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_5_i_clk clknet_4_2_0_i_clk VGND VGND VPWR VPWR clknet_leaf_5_i_clk sky130_fd_sc_hd__clkbuf_16
X_14776_ clknet_leaf_76_i_clk _00321_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11988_ _05092_ _05105_ _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13727_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06602_
+ _06562_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__o21ai_1
X_10939_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04177_ VGND
+ VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13658_ _06200_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06545_
+ _06546_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12609_ _05621_ _05637_ _05629_ _05597_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__or4bb_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13589_ _06472_ _06474_ _06481_ _06480_ _06471_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__o311a_1
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15328_ clknet_leaf_19_i_clk _00873_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15259_ clknet_leaf_3_i_clk _00804_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09820_ _03211_ _03212_ _02850_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__mux2_1
X_09751_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03142_ _03154_
+ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__o21ai_1
X_08702_ _02222_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09682_ _03072_ _03081_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08633_ _02158_ _02160_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[15\] _02099_ VGND VGND VPWR
+ VPWR _02100_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07515_ _01229_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08495_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[8\] _02036_ VGND VGND VPWR
+ VPWR _02037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07446_ _01177_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07377_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _01051_ _01052_
+ _01116_ _01057_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09116_ _02585_ _02583_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_134_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09047_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _02527_ VGND
+ VGND VPWR VPWR _02528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold450 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND VGND VPWR
+ VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold483 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _06297_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
X_09949_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03315_ _03205_
+ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__o21a_1
X_12960_ _05843_ _05936_ _05937_ _05938_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__o211a_1
X_11911_ _05036_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__nand2_1
X_12891_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR _05881_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ clknet_leaf_44_i_clk _00175_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _04930_ VGND
+ VGND VPWR VPWR _04976_ sky130_fd_sc_hd__xnor2_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ clknet_leaf_41_i_clk _00107_ VGND VGND VPWR VPWR diff2\[5\] sky130_fd_sc_hd__dfxtp_1
X_11773_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13512_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _06352_ VGND
+ VGND VPWR VPWR _06418_ sky130_fd_sc_hd__xnor2_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _03995_ net186 _04003_ _04004_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ clknet_leaf_4_i_clk _00038_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13443_ _06345_ _06350_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10655_ _03910_ _03915_ _03925_ _03937_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13374_ _06295_ net610 _06216_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__a21o_1
X_10586_ _03882_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15113_ clknet_leaf_112_i_clk _00658_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12325_ _05392_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15044_ clknet_leaf_104_i_clk _00589_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12256_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _05291_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__o21ai_1
X_11207_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _04398_ VGND VGND
+ VPWR VPWR _04420_ sky130_fd_sc_hd__and4_1
X_12187_ _05241_ _05246_ _05247_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11138_ _03976_ _04368_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__and2_1
X_11069_ _04305_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14828_ clknet_leaf_77_i_clk _00373_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14759_ clknet_leaf_64_i_clk _00304_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07300_ _01046_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__buf_2
X_08280_ _01748_ _01850_ _01851_ _01472_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07231_ _00994_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_106_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_106_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09803_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] _03193_
+ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07995_ _01463_ net638 _01460_ _01596_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09734_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _03140_ sky130_fd_sc_hd__or2_1
X_09665_ _02746_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _03075_
+ _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__a22o_1
X_08616_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR VPWR
+ _02146_ sky130_fd_sc_hd__inv_2
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08547_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\] _02084_ VGND VGND VPWR
+ VPWR _02085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08478_ _02021_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07429_ _01161_ _01162_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10440_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03651_ _03745_
+ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_123_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10371_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03650_ VGND VGND VPWR
+ VPWR _03690_ sky130_fd_sc_hd__o31a_1
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12110_ _05130_ _05202_ _05204_ _05080_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__o211a_1
X_13090_ _06028_ _06052_ _06050_ net112 _05860_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a41o_1
XFILLER_0_103_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12041_ _04829_ _05144_ _05145_ _05129_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__a31o_1
Xhold280 diff2\[3\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND VPWR
+ VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_70_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13992_ _06555_ _06831_ _06832_ _06747_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__o211a_1
X_12943_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05923_
+ _05842_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12874_ _05854_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _05865_ _05866_ _05751_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _04951_ _04960_ _04961_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__o21a_1
X_14613_ clknet_leaf_42_i_clk _00158_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14544_ clknet_leaf_33_i_clk _00090_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
X_11756_ _04773_ net443 _04898_ _04899_ _04788_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o221a_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10707_ _03992_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14475_ clknet_leaf_7_i_clk _00021_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_1
X_11687_ _04832_ _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13426_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _06342_
+ _06343_ _06285_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__o221a_1
X_10638_ _03535_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13357_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06282_
+ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__and2_1
X_10569_ _03621_ net510 VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12308_ _05374_ _05378_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_23_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13288_ _05928_ _06218_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15027_ clknet_leaf_97_i_clk _00572_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12239_ _05317_ _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_38_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07780_ net189 _01345_ _01336_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 in_alpha[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
X_09450_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__or4_2
XFILLER_0_59_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08401_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[15\] _01946_ _01882_
+ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09381_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _02817_
+ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08332_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[5\] _01894_ VGND VGND
+ VPWR VPWR _01895_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08263_ net42 net24 VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08194_ _01565_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07978_ _01565_ _01567_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__o21ai_1
X_09717_ _03122_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09648_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03060_ VGND
+ VGND VPWR VPWR _03061_ sky130_fd_sc_hd__and2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _02986_ VGND
+ VGND VPWR VPWR _02999_ sky130_fd_sc_hd__or2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _04769_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _04762_ _04772_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__o211a_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _05619_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11541_ _04712_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14260_ _06910_ net587 _06678_ _07060_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11472_ _04651_ _04653_ _04655_ _04374_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13211_ _06138_ _06141_ _06150_ _06155_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__and4_1
X_10423_ _03623_ _03736_ _03737_ _03515_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__o211a_1
X_14191_ _06875_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _06904_
+ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13142_ _05854_ net270 _05847_ _06099_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10354_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _03674_ VGND
+ VGND VPWR VPWR _03675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13073_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _06003_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__o21ai_1
X_10285_ _03607_ net124 _03568_ _03618_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__o211a_1
X_12024_ net153 _05132_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__or2_1
X_13975_ _06816_ _06817_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12926_ _05871_ net627 _05908_ _05909_ _05910_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _05843_ net176 _05847_ _05852_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__o211a_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _04862_ _04945_ _04946_ _04739_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12788_ _05795_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__xor2_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11739_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _04864_ _04794_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__o31a_1
X_14527_ clknet_leaf_42_i_clk _00073_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14458_ clknet_leaf_40_i_clk _00004_ VGND VGND VPWR VPWR r_i_alpha1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13409_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _06326_ VGND
+ VGND VPWR VPWR _06328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14389_ _07169_ _07170_ _07171_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08950_ _02439_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07901_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\] _01498_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\]
+ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__o21a_1
X_08881_ _02314_ _02379_ _02380_ _02260_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__o211a_1
X_07832_ net203 _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__or2_1
X_07763_ net10 _01405_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09502_ _02923_ _02928_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07694_ _01359_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09433_ _02865_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _02807_ _02808_ _02409_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08315_ _01879_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_4
X_09295_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08246_ _01662_ _01820_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08177_ _01529_ net454 _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10070_ _03431_ _03432_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__and2b_1
X_13760_ _01474_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__clkbuf_4
X_10972_ _04011_ net282 _04003_ _04218_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__o211a_1
X_12711_ _05359_ _05712_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13691_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND VPWR
+ VPWR _06572_ sky130_fd_sc_hd__a21oi_1
X_12642_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05641_ VGND
+ VGND VPWR VPWR _05667_ sky130_fd_sc_hd__or2_1
X_15430_ clknet_leaf_8_i_clk _00975_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15361_ clknet_leaf_21_i_clk _00906_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_12573_ _05488_ _05604_ _05605_ _05343_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11524_ _04468_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__and2_1
X_14312_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _07042_ VGND
+ VGND VPWR VPWR _07105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15292_ clknet_leaf_17_i_clk _00837_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14243_ _07044_ _07045_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__and2_1
X_11455_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _04639_ VGND
+ VGND VPWR VPWR _04640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10406_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03721_ VGND
+ VGND VPWR VPWR _03722_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14174_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _06985_
+ _01862_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04565_ VGND
+ VGND VPWR VPWR _04580_ sky130_fd_sc_hd__or2_1
X_13125_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06083_ VGND
+ VGND VPWR VPWR _06084_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10337_ _03642_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__nand2_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _05998_ _06023_ _06024_ _05938_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__o211a_1
X_10268_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _03609_
+ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__or2_1
X_12007_ _05123_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_1
X_10199_ _03105_ _03538_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__nor2_1
X_13958_ _06501_ _06802_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12909_ _05566_ _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13889_ _06556_ _06741_ _06742_ _06459_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08100_ _01669_ _01693_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09080_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08031_ _01627_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__xnor2_1
Xinput40 in_y[10] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 in_y[4] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09982_ _03306_ _03310_ _03335_ _03336_ _03346_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__o2111a_1
X_08933_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02423_ VGND
+ VGND VPWR VPWR _02424_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08864_ _01958_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__or2_1
X_07815_ _01444_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
X_08795_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _01876_ _02306_
+ _02307_ _02309_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07746_ _01395_ _01396_ net194 _01345_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__a2bb2o_1
X_07677_ _01334_ _01341_ net18 VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09416_ _02845_ _02852_ _02747_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09347_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02788_
+ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09278_ _02733_ _02735_ _02312_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08229_ _01625_ _01646_ _01809_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11240_ _04447_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _04448_ sky130_fd_sc_hd__nor2_1
X_11171_ _04378_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10122_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03478_ VGND
+ VGND VPWR VPWR _03479_ sky130_fd_sc_hd__xor2_1
X_14930_ clknet_leaf_81_i_clk _00475_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_10053_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03410_ VGND
+ VGND VPWR VPWR _03418_ sky130_fd_sc_hd__nand2_1
X_14861_ clknet_leaf_85_i_clk _00406_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13812_ _06673_ _06674_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__xor2_1
X_14792_ clknet_leaf_66_i_clk _00337_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10955_ _04202_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__or2_1
X_13743_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06611_
+ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10886_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _04142_ sky130_fd_sc_hd__inv_2
X_13674_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _06557_
+ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15413_ clknet_leaf_26_i_clk _00958_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12625_ _01252_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__buf_2
XFILLER_0_156_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12556_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05589_ VGND
+ VGND VPWR VPWR _05590_ sky130_fd_sc_hd__and2_1
X_15344_ clknet_leaf_48_i_clk _00889_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11507_ _04685_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12487_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _05531_
+ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15275_ clknet_leaf_17_i_clk _00820_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold109 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _04624_ _04615_ _04612_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__a21o_1
X_14226_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _07021_ VGND
+ VGND VPWR VPWR _07031_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14157_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _06967_
+ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11369_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04414_ _04564_
+ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__o21ai_4
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _05854_ net294 _05847_ _06068_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__o211a_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__or2_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _06003_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07600_ r_i_alpha1\[6\] _01285_ _01276_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__mux2_1
X_08580_ _02101_ _02107_ _02114_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07531_ net73 net348 _01234_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07462_ _01044_ net374 _01189_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09201_ _02664_ _02666_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07393_ _01129_ _01130_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09132_ _02312_ _02602_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09063_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02541_ VGND
+ VGND VPWR VPWR _02542_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08014_ _01598_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09965_ _03314_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__a21oi_1
X_08916_ net531 _02405_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__nand2_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03260_ _03207_
+ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__o41a_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02351_
+ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08778_ _02282_ _02285_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__a21oi_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ net18 _01341_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ _03958_ _03961_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12410_ _05463_ _05465_ _05469_ _05222_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13390_ _06307_ _06309_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12341_ _05397_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15060_ clknet_leaf_112_i_clk _00605_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12272_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14011_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06837_ VGND
+ VGND VPWR VPWR _06849_ sky130_fd_sc_hd__or2_1
X_11223_ _04414_ _04432_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11154_ net128 _04379_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__or2_1
X_10105_ _03024_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__and2_1
X_11085_ _04047_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04320_
+ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a22o_1
X_14913_ clknet_leaf_81_i_clk _00458_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_10036_ _03396_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__or2_1
X_14844_ clknet_leaf_86_i_clk _00389_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14775_ clknet_leaf_76_i_clk _00320_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_11987_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _05081_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13726_ _06293_ _06599_ _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__o21a_1
X_10938_ _03801_ _04188_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10869_ _04048_ _04125_ _04126_ _04063_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__o211a_1
X_13657_ _06518_ _06544_ _06540_ _06541_ _06199_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__a41oi_1
XFILLER_0_128_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12608_ _05603_ _05608_ _05609_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__nand3_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13588_ _01765_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15327_ clknet_leaf_17_i_clk _00872_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_12539_ _05570_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15258_ clknet_leaf_10_i_clk _00803_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14209_ _01253_ _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__and2_1
X_15189_ clknet_leaf_124_i_clk _00734_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09750_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03144_ _03142_
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND VPWR VPWR
+ _03154_ sky130_fd_sc_hd__a22o_1
X_08701_ _02213_ _02223_ _02211_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__o21ai_1
X_09681_ _03051_ _03061_ _03062_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_146_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08632_ _02158_ _02160_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08563_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\]
+ _02083_ _01881_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07514_ net416 _01228_ _01013_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08494_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\] _02035_ VGND VGND VPWR
+ VPWR _02036_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07445_ net76 _01176_ _01013_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07376_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _01108_ VGND
+ VGND VPWR VPWR _01116_ sky130_fd_sc_hd__xor2_1
X_09115_ _02152_ _02587_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09046_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _02526_ VGND
+ VGND VPWR VPWR _02527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold440 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold451 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND VGND VPWR
+ VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _00841_ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
X_09948_ _03184_ _03321_ _03322_ _03292_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__o211a_1
X_09879_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03261_
+ _03186_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__o21ai_1
X_11910_ _05033_ _05035_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__nand2_1
X_12890_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _05862_ _05878_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a31o_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _04966_ _04971_ _04967_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__a21boi_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _04913_ _04795_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__mux2_1
X_14560_ clknet_leaf_39_i_clk _00106_ VGND VGND VPWR VPWR diff2\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] _03999_
+ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__or2_1
X_13511_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06352_ _06414_
+ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__a21o_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ clknet_leaf_4_i_clk _00037_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13442_ _06329_ _06338_ _06339_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__and3_1
X_10654_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03945_ VGND
+ VGND VPWR VPWR _03946_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13373_ _06295_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _06296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10585_ _03680_ _03881_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15112_ clknet_leaf_113_i_clk net343 VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12324_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _05393_ VGND
+ VGND VPWR VPWR _05394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15043_ clknet_leaf_104_i_clk _00588_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12255_ _05308_ _05319_ _05320_ _05326_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11206_ _04390_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _04418_ _04419_ _04360_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__o221a_1
X_12186_ _05255_ _05270_ _05265_ _05271_ _05264_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__o32a_1
XFILLER_0_102_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11137_ _04047_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04366_
+ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__a22o_1
X_11068_ _04291_ _04297_ _04295_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__o21ai_1
X_10019_ _03383_ _03379_ _03386_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14827_ clknet_leaf_77_i_clk _00372_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14758_ clknet_leaf_64_i_clk _00303_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ _06586_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14689_ clknet_leaf_57_i_clk _00234_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_07230_ net365 _00991_ _00993_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09802_ net136 _03189_ _03017_ _03197_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07994_ _01556_ _01592_ _01594_ _01595_ _01485_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09733_ _03133_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__xnor2_1
X_09664_ _03061_ _03067_ _03074_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__o31a_1
X_08615_ _01961_ _02140_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__nor2_1
X_09595_ _02844_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03011_
+ _03012_ _03013_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__o221a_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _01881_ _02083_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08477_ _01981_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07428_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _01160_ VGND
+ VGND VPWR VPWR _01162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07359_ _01099_ _01100_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__and2_1
X_10370_ _03679_ _03689_ _02132_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09029_ _02497_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_i_clk clknet_4_2_0_i_clk VGND VGND VPWR VPWR clknet_leaf_4_i_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ _05144_ _05145_ _04829_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold270 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold281 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] VGND VGND
+ VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
X_13991_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND
+ VGND VPWR VPWR _06832_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12942_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05923_
+ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _05859_ _05864_ _05842_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a21o_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ clknet_leaf_45_i_clk _00157_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _01794_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__buf_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ clknet_leaf_39_i_clk _00089_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_11755_ _04886_ _04889_ _04897_ _04755_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10706_ _03642_ _02310_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14474_ clknet_leaf_5_i_clk _00020_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
X_11686_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _04835_ VGND
+ VGND VPWR VPWR _04836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13425_ _06340_ _06341_ _06205_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__o21ai_1
X_10637_ _03929_ _03930_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ _03605_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10568_ _03860_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__xor2_1
X_13356_ _05928_ _06279_ _06281_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12307_ _05374_ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10499_ _03805_ _03806_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__and2_1
X_13287_ _06204_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__clkbuf_4
X_15026_ clknet_leaf_97_i_clk _00571_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12238_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05291_ VGND
+ VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nand2_1
X_12169_ _05246_ _05252_ _05255_ _05128_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 in_alpha[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08400_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[15\] _01947_ _01882_
+ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09380_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _02819_
+ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08331_ _01892_ _01893_ _01882_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08262_ _01465_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\] _01836_ _01837_
+ _01661_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08193_ _01553_ _01570_ _01569_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07977_ net31 net49 VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__nand2_1
X_09716_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03121_ VGND
+ VGND VPWR VPWR _03123_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09647_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03059_ VGND
+ VGND VPWR VPWR _03060_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09578_ _02844_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _02997_
+ _02998_ _02827_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__o221a_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08529_ _01865_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02067_
+ _02068_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11540_ _04714_ _04716_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11471_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _04639_ _04654_
+ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13210_ _06158_ _06159_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__and2b_1
X_10422_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _03737_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14190_ _06875_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _06999_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13141_ _05855_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nand2_1
X_10353_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13072_ _06025_ _06032_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__or2_1
X_10284_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _03609_
+ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__or2_1
X_12023_ _05130_ net257 _04979_ _05134_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__o211a_1
X_13974_ _06804_ _06811_ _06809_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__a21o_1
X_12925_ _04538_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__clkbuf_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05845_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _04765_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _04946_ sky130_fd_sc_hd__or2_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _05786_ _05790_ _05787_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__o21bai_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_105_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_105_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ clknet_leaf_46_i_clk _00072_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11738_ _04868_ _04875_ _04876_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14457_ clknet_leaf_41_i_clk _00003_ VGND VGND VPWR VPWR r_i_alpha1\[7\] sky130_fd_sc_hd__dfxtp_1
X_11669_ _04773_ net606 _04821_ _04822_ _04788_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13408_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _06326_ VGND
+ VGND VPWR VPWR _06327_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14388_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _07156_ VGND
+ VGND VPWR VPWR _07171_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13339_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _06266_ _06267_ _06197_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15009_ clknet_leaf_108_i_clk _00554_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_07900_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[10\] _01510_
+ _01511_ _01513_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__o221a_1
X_08880_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07831_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in VGND VGND VPWR VPWR _01457_
+ sky130_fd_sc_hd__clkbuf_4
X_07762_ net10 _01405_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__or2_1
X_09501_ _02923_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__or2_1
X_07693_ net337 _01357_ _01358_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09432_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02864_ VGND
+ VGND VPWR VPWR _02866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09363_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _02800_
+ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08314_ _01549_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__inv_2
X_09294_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _02750_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08245_ _01455_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08176_ _01765_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_84_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_99_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_99_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10971_ _04216_ _04217_ _04012_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__o21ai_1
X_12710_ _05724_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13690_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND VPWR
+ VPWR _06571_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12641_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05641_ VGND
+ VGND VPWR VPWR _05666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15360_ clknet_leaf_20_i_clk _00905_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12572_ _05492_ net498 VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14311_ _07089_ _07103_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__nor2_1
X_11523_ _04378_ _04700_ _04701_ _04702_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__a31o_1
X_15291_ clknet_leaf_17_i_clk _00836_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_37_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14242_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _07023_ VGND
+ VGND VPWR VPWR _07045_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11454_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04638_ VGND
+ VGND VPWR VPWR _04639_ sky130_fd_sc_hd__xor2_2
XFILLER_0_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10405_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03720_ VGND
+ VGND VPWR VPWR _03721_ sky130_fd_sc_hd__xnor2_1
X_11385_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04565_ VGND
+ VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nand2_1
X_14173_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _06985_
+ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13124_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05878_ VGND VGND
+ VPWR VPWR _06083_ sky130_fd_sc_hd__o31a_1
X_10336_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _03660_
+ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__xnor2_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _03608_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__buf_2
X_13055_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND
+ VGND VPWR VPWR _06024_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12006_ _04850_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__and2_1
X_10198_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03547_ VGND
+ VGND VPWR VPWR _03548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13957_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _06801_ _06553_
+ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__mux2_1
X_12908_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _05884_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13888_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _06742_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12839_ _05490_ _02310_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__and2_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14509_ clknet_leaf_31_i_clk _00055_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08030_ _01612_ _01620_ _01628_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 in_x[1] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
Xinput41 in_y[11] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput52 in_y[5] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09981_ _03335_ _03337_ _03346_ _03351_ _03345_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__a32o_1
X_08932_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _02422_ VGND
+ VGND VPWR VPWR _02423_ sky130_fd_sc_hd__xnor2_1
X_08863_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02349_
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07814_ net426 _01443_ _01411_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__mux2_1
X_08794_ _02308_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__clkbuf_4
X_07745_ net5 _01393_ _01338_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__o21ai_1
X_07676_ _01334_ net18 _01341_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09415_ net440 _02846_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09346_ _02754_ net357 _02749_ _02793_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09277_ _02733_ _02735_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08228_ _01599_ _01643_ _01791_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08159_ _01748_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11170_ _04377_ net290 _04387_ _04389_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10121_ _03205_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10052_ _03191_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03416_
+ _03417_ _03258_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14860_ clknet_leaf_86_i_clk _00405_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13811_ _06663_ _06665_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__nand2_1
X_14791_ clknet_leaf_68_i_clk _00336_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13742_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06600_ VGND VGND
+ VPWR VPWR _06615_ sky130_fd_sc_hd__and4_1
X_10954_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04177_ VGND
+ VGND VPWR VPWR _04203_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13673_ _06556_ net212 _06485_ _06558_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__o211a_1
X_10885_ _04048_ _04140_ _04141_ _04063_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15412_ clknet_leaf_28_i_clk _00957_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_12624_ _05632_ _05650_ _05651_ _05343_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15343_ clknet_leaf_38_i_clk _00888_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12555_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05588_ VGND
+ VGND VPWR VPWR _05589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11506_ _04686_ _04680_ _04674_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15274_ clknet_leaf_13_i_clk _00819_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12486_ _05530_ _05528_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14225_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _07023_ VGND
+ VGND VPWR VPWR _07030_ sky130_fd_sc_hd__nand2_1
X_11437_ _04233_ _04610_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14156_ _06910_ net236 _06678_ _06971_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__o211a_1
X_11368_ _04061_ _04543_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__or2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _06066_ _06067_ _05855_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _03644_ _03645_ _03280_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__mux2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__nand2_1
X_11299_ _04413_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__and2_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05982_ VGND
+ VGND VPWR VPWR _06009_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14989_ clknet_leaf_107_i_clk _00534_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_135_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07530_ _01237_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07461_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _01159_ _01187_
+ _01188_ _01059_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09200_ _02655_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07392_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _01119_ VGND
+ VGND VPWR VPWR _01130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09131_ _02596_ _02589_ _02601_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09062_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _02540_ VGND
+ VGND VPWR VPWR _02541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08013_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09964_ _03318_ _03325_ _03326_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__o21a_1
X_08915_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _02409_ sky130_fd_sc_hd__clkbuf_4
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _03271_ _03264_ _03253_ _03266_ _02850_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__o41a_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _02348_ _02350_ _02344_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__mux2_1
X_08777_ _02282_ _02285_ _02275_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__o21a_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ net224 _01333_ _01382_ _01383_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__o22a_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07659_ _01332_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10670_ _03957_ _03955_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09329_ _02409_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _02776_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12340_ _05407_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12271_ _05140_ net272 _05141_ _05346_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__o211a_1
X_14010_ _06555_ _06847_ _06848_ _06747_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__o211a_1
X_11222_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04420_ _04414_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__a31o_1
X_11153_ _04377_ net157 _04219_ _04380_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10104_ _03182_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _03461_
+ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a22o_1
X_11084_ _04319_ _04309_ _04312_ _03993_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__a31oi_1
X_14912_ clknet_leaf_81_i_clk _00457_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10035_ _03364_ _03374_ _03397_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__o31a_1
X_14843_ clknet_leaf_85_i_clk _00388_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14774_ clknet_leaf_52_i_clk _00319_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11986_ _05095_ _05099_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13725_ _06292_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__nand2_1
X_10937_ _04177_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13656_ _06518_ _06540_ _06541_ _06544_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10868_ _04010_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _04126_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ _05619_ _05628_ _05634_ _05621_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__o221a_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ _06201_ _06483_ _06484_ _06459_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__o211a_1
X_10799_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _04064_ sky130_fd_sc_hd__inv_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15326_ clknet_leaf_17_i_clk _00871_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12538_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _05573_ VGND
+ VGND VPWR VPWR _05574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15257_ clknet_leaf_10_i_clk _00802_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12469_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _05504_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__or3_1
X_14208_ _06903_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _07013_
+ _07014_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15188_ clknet_leaf_124_i_clk _00733_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14139_ _06646_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _06946_ _06956_
+ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__o41a_1
XFILLER_0_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08700_ _02194_ _02214_ _02216_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a21oi_1
X_09680_ _02891_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08631_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[4\] _02159_ VGND VGND VPWR
+ VPWR _02160_ sky130_fd_sc_hd__xnor2_1
X_08562_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _02097_
+ _02098_ _02055_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__o221a_1
X_07513_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _01026_ _01226_
+ _01227_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08493_ _01880_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07444_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ _01010_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07375_ _01019_ _01114_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09114_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _02586_ VGND
+ VGND VPWR VPWR _02587_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09045_ _02343_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold430 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _00778_ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold463 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold474 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\] VGND VGND VPWR VPWR
+ net613 sky130_fd_sc_hd__dlygate4sd3_1
X_09947_ _03290_ net614 VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__or2_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _03261_
+ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08829_ _01958_ _02335_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _04974_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04904_ _04794_
+ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _06409_ _06416_ _04961_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__o21a_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _03619_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14490_ clknet_leaf_4_i_clk _00036_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13441_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ _06351_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__o21ai_1
X_10653_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03941_ _03944_
+ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13372_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND VGND
+ VPWR VPWR _06295_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10584_ _03680_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15111_ clknet_leaf_112_i_clk _00656_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12323_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ _05375_ _05163_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15042_ clknet_leaf_104_i_clk _00587_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_12254_ _05330_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11205_ _04417_ _04415_ _04416_ _04396_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__a31o_1
X_12185_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05254_ _05263_
+ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11136_ _04365_ _04361_ _04362_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__o31a_1
X_11067_ _04303_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__nand2_1
X_10018_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03385_ VGND
+ VGND VPWR VPWR _03386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14826_ clknet_leaf_110_i_clk _00371_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14757_ clknet_leaf_65_i_clk _00302_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11969_ _04771_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05089_
+ _05090_ _04965_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__o221a_1
X_13708_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _06586_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14688_ clknet_leaf_55_i_clk _00233_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13639_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _06514_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15309_ clknet_leaf_23_i_clk _00854_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09801_ _03195_ _03196_ _03191_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07993_ _01589_ _01593_ _01572_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__a21o_1
X_09732_ _03123_ _03134_ _03136_ _03094_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__a221o_2
X_09663_ _03061_ _03067_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__o21ai_2
X_08614_ _01876_ net310 _01945_ _02144_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09594_ _02308_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\]
+ _02056_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08476_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02019_ _01868_
+ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07427_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _01160_ VGND
+ VGND VPWR VPWR _01161_ sky130_fd_sc_hd__or2_1
X_07358_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _01082_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _01010_
+ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09028_ _02319_ _02508_ _02509_ _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold260 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\] VGND VGND VPWR VPWR
+ net410 sky130_fd_sc_hd__dlygate4sd3_1
X_13990_ _06829_ _06830_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__xnor2_1
X_12941_ _05921_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2b_1
X_12872_ _05859_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__nor2_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ clknet_leaf_46_i_clk _00156_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _04958_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__nor2_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ clknet_leaf_38_i_clk _00088_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _04886_ _04889_ _04897_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__a21oi_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10705_ net535 _03625_ _03990_ _03991_ _03814_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__o221a_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ clknet_leaf_5_i_clk _00019_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11685_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04834_ VGND
+ VGND VPWR VPWR _04835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13424_ _06340_ _06341_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__and2_1
X_10636_ _03927_ _03928_ _03925_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13355_ _05927_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__nand2_1
X_10567_ _03865_ _03866_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _05377_ VGND
+ VGND VPWR VPWR _05378_ sky130_fd_sc_hd__xnor2_1
X_13286_ _06210_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _06221_ _06222_ _06197_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__o221a_1
X_10498_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03796_ VGND
+ VGND VPWR VPWR _03806_ sky130_fd_sc_hd__or2_1
X_15025_ clknet_leaf_97_i_clk _00570_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_12237_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05279_ VGND
+ VGND VPWR VPWR _05317_ sky130_fd_sc_hd__or2_1
X_12168_ _05246_ _05252_ _05255_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__a21o_1
X_11119_ _04132_ _04338_ _04336_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__a22o_1
X_12099_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05194_
+ _01250_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__o21ai_1
Xinput6 in_alpha[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_0_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14809_ clknet_leaf_67_i_clk _00354_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND VPWR VPWR _01893_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08261_ _01330_ _01712_ _01529_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08192_ _01539_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\] _01778_ _01779_
+ _01661_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07976_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_2
X_09715_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03121_ VGND
+ VGND VPWR VPWR _03122_ sky130_fd_sc_hd__nand2_1
X_09646_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _03048_ _02770_
+ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _02993_ _02989_ _02996_ _02761_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__a31o_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08528_ _02061_ _02066_ _01868_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08459_ _02002_ _02003_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11470_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _04641_ _04639_
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR VPWR
+ _04654_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10421_ _03734_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13140_ _06093_ _06097_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10352_ _03626_ net569 _03672_ _03673_ _03633_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13071_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06003_ VGND
+ VGND VPWR VPWR _06037_ sky130_fd_sc_hd__xnor2_2
X_10283_ _03607_ net126 _03568_ _03617_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12022_ net149 _05132_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__or2_1
X_13973_ _06814_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__and2b_1
X_12924_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _05907_
+ _05845_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__o21ai_1
X_12855_ _05843_ net167 _05847_ _05851_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__o211a_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _04941_ _04944_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _05793_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__nor2_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ clknet_leaf_47_i_clk _00071_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.i_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11737_ _04863_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__and2_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_899 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14456_ clknet_leaf_41_i_clk _00002_ VGND VGND VPWR VPWR r_i_alpha1\[6\] sky130_fd_sc_hd__dfxtp_1
X_11668_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04820_
+ _04755_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13407_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06325_ VGND
+ VGND VPWR VPWR _06326_ sky130_fd_sc_hd__xor2_1
X_10619_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03913_ VGND
+ VGND VPWR VPWR _03914_ sky130_fd_sc_hd__xor2_2
XFILLER_0_4_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14387_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ _07156_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__o41a_1
X_11599_ _04757_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13338_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06265_
+ _06232_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13269_ _06205_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ clknet_leaf_103_i_clk _00553_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07830_ _01455_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__buf_4
X_07761_ _01405_ _01407_ net262 _01345_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__a2bb2o_1
X_09500_ _02907_ _02898_ _02914_ _02927_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07692_ _00992_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02864_ VGND
+ VGND VPWR VPWR _02865_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_3_i_clk clknet_4_2_0_i_clk VGND VGND VPWR VPWR clknet_leaf_3_i_clk sky130_fd_sc_hd__clkbuf_16
X_09362_ _02806_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08313_ _01876_ net307 _01823_ _01878_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09293_ _01455_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08244_ _01717_ net475 _01635_ _01822_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08175_ _01251_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07959_ net49 net31 VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10970_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__nor2_1
X_09629_ _02745_ _03042_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12640_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05664_
+ _05665_ _05544_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12571_ _05597_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14310_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _07042_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11522_ _04375_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND
+ VGND VPWR VPWR _04702_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15290_ clknet_leaf_16_i_clk _00835_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14241_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _07023_ VGND
+ VGND VPWR VPWR _07044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11453_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] net652 _04412_
+ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10404_ net117 _03719_ _03280_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14172_ _06983_ _06984_ _06934_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__mux2_1
X_11384_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _04565_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13123_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _06082_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10335_ _03657_ _03659_ _03651_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__mux2_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _06021_ _06022_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__xnor2_1
X_10266_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _03608_ sky130_fd_sc_hd__buf_2
X_12005_ _04754_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05120_
+ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__a22o_1
X_10197_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03546_ VGND
+ VGND VPWR VPWR _03547_ sky130_fd_sc_hd__xor2_2
X_13956_ _06799_ _06800_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__xnor2_1
X_12907_ _05843_ _05893_ _05894_ _05675_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__o211a_1
X_13887_ _06736_ _06740_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__xor2_1
X_12838_ _05632_ _05838_ _05839_ _05675_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__o211a_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12769_ _05732_ _05761_ _05752_ _05774_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14508_ clknet_leaf_31_i_clk _00054_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 in_alpha[9] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
X_14439_ _07208_ _07210_ _07213_ _06926_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__a31o_1
Xinput31 in_x[2] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
Xinput42 in_y[12] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 in_y[6] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09980_ _03347_ _03344_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08931_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _02422_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08862_ _01959_ _02363_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__nand2_1
X_07813_ net8 _01441_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__xor2_1
X_08793_ _01252_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__clkbuf_4
X_07744_ net5 _01393_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__and2_1
X_07675_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_4
X_09414_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09345_ _02755_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09276_ _02717_ _02721_ _02730_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__o31a_1
XFILLER_0_74_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08227_ _01465_ net511 _01807_ _01808_ _01661_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08158_ _01746_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__or2_2
XFILLER_0_101_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08089_ _01681_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10120_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__or4_2
XFILLER_0_101_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10051_ _03414_ _03415_ _03186_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_104_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_104_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13810_ _06671_ _06672_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__and2_1
X_14790_ clknet_leaf_66_i_clk _00335_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_119_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13741_ _06565_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _06613_ _06614_ _06526_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__o221a_1
X_10953_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04177_ VGND
+ VGND VPWR VPWR _04202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13672_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _06557_
+ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10884_ _04010_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _04141_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12623_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND
+ VGND VPWR VPWR _05651_ sky130_fd_sc_hd__or2_1
X_15411_ clknet_leaf_24_i_clk _00956_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_156_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15342_ clknet_leaf_38_i_clk _00887_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12554_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05526_ VGND VGND
+ VPWR VPWR _05588_ sky130_fd_sc_hd__o31a_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11505_ _04676_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15273_ clknet_leaf_11_i_clk _00818_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12485_ _05522_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14224_ _07024_ _07026_ _07022_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11436_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14155_ _06966_ _06969_ _06970_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__o21ai_1
X_11367_ _04529_ _04535_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ _06060_ _06065_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__and2_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03634_
+ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__nand2_1
X_14086_ _06910_ net245 _06678_ _06912_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__o211a_1
X_11298_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ _04481_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__or3_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _05998_ _06007_ _06008_ _05938_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__o211a_1
X_10249_ _03574_ _03577_ _03592_ _03572_ _03390_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14988_ clknet_leaf_104_i_clk _00533_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13939_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06784_ VGND
+ VGND VPWR VPWR _06785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07460_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _01122_ _01063_
+ _01047_ _01057_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_83_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07391_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _01119_ VGND
+ VGND VPWR VPWR _01129_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09130_ _02596_ _02589_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09061_ _02344_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_98_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08012_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__buf_2
XFILLER_0_142_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_i_clk clknet_4_8_0_i_clk VGND VGND VPWR VPWR clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09963_ _03320_ _03327_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__and2_1
X_08914_ _02387_ net440 _02407_ _02408_ _02309_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__o221a_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _03184_ _03274_ _03275_ _03058_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__o211a_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _02349_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__inv_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08776_ _02257_ _02271_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__and3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _01338_ _01341_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07658_ _01059_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07589_ r_i_alpha1\[4\] _01275_ _01276_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09328_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _02777_
+ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09259_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _02704_ _02719_
+ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12270_ _05344_ _05345_ _05142_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_133_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11221_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04427_
+ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__or2_1
X_11152_ net143 _04379_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10103_ _03458_ _03460_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__o21a_1
X_11083_ _04309_ _04312_ _04319_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a21o_1
X_14911_ clknet_leaf_81_i_clk _00456_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10034_ _03377_ _03397_ _03399_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__o22a_1
X_14842_ clknet_leaf_85_i_clk _00387_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11985_ _05102_ _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__nor2_1
X_14773_ clknet_leaf_53_i_clk _00318_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10936_ _04023_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04186_
+ _04187_ _04059_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__o221a_1
X_13724_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _06593_
+ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10867_ _04123_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__xnor2_1
X_13655_ _06542_ _06543_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _05627_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13586_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND
+ VGND VPWR VPWR _06484_ sky130_fd_sc_hd__or2_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ _04048_ _04060_ _04062_ _04063_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__o211a_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12537_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05572_ VGND
+ VGND VPWR VPWR _05573_ sky130_fd_sc_hd__xnor2_1
X_15325_ clknet_leaf_18_i_clk _00870_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12468_ _05500_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _05514_ _05515_ _05391_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__o221a_1
X_15256_ clknet_leaf_5_i_clk _00801_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11419_ _04444_ net591 VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__or2_1
X_14207_ _07010_ _07012_ _01861_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__o21a_1
X_15187_ clknet_leaf_123_i_clk _00732_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12399_ _05434_ _05448_ _05453_ _05456_ _05449_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_22_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14138_ _06647_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _06951_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14069_ _06893_ _06895_ _06898_ _06569_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__a31o_1
X_08630_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\] _01879_ VGND VGND VPWR VPWR
+ _02159_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08561_ _02095_ _02096_ _01866_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07512_ _01010_ _01172_ _01037_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__a2bb2o_1
X_08492_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[6\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\]
+ _01992_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__or4_4
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07443_ _01095_ net306 _01174_ _01175_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07374_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _01105_ VGND
+ VGND VPWR VPWR _01114_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09113_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ _02341_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09044_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _02504_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold420 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold431 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold442 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND VPWR
+ VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR
+ VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold464 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND VGND VPWR
+ VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold497 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09946_ _03314_ _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__xor2_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _03253_ _03259_ _03260_ _02850_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__o22a_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08828_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND VPWR
+ VPWR _02335_ sky130_fd_sc_hd__and3_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _02275_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__nand2_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _04769_ net389 _04762_ _04912_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__o211a_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _03995_ net277 _03620_ _04002_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__o211a_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _06211_ net593 _06354_ _06355_ _06285_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__o221a_1
X_10652_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13371_ _06202_ _06291_ _06294_ _06110_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__o211a_1
X_10583_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03880_ VGND
+ VGND VPWR VPWR _03881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12322_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _05392_ sky130_fd_sc_hd__inv_2
X_15110_ clknet_leaf_112_i_clk _00655_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15041_ clknet_leaf_103_i_clk _00586_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12253_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05291_ VGND
+ VGND VPWR VPWR _05331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11204_ _04415_ _04416_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12184_ _05239_ _05269_ _05247_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__o21ai_1
X_11135_ _04361_ _04362_ _04365_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11066_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04302_ VGND
+ VGND VPWR VPWR _04304_ sky130_fd_sc_hd__or2_1
X_10017_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03384_ VGND
+ VGND VPWR VPWR _03385_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14825_ clknet_leaf_110_i_clk _00370_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14756_ clknet_leaf_64_i_clk _00301_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_4
X_11968_ _05087_ _05088_ _04786_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13707_ _06565_ net590 _06583_ _06585_ _06526_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__o221a_1
X_10919_ _04023_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04171_
+ _04172_ _04059_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__o221a_1
X_11899_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05026_ VGND
+ VGND VPWR VPWR _05027_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14687_ clknet_leaf_54_i_clk _00232_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13638_ _06527_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13569_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND
+ VGND VPWR VPWR _06469_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15308_ clknet_leaf_22_i_clk _00853_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15239_ clknet_leaf_11_i_clk _00784_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09800_ _03193_ _03194_ _02851_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__a21oi_1
X_07992_ _01589_ _01593_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09731_ _03114_ _03135_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09662_ _03072_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__and2_2
XFILLER_0_97_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08613_ _02142_ _02143_ _01877_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__o21ai_1
X_09593_ _03000_ _03009_ _03010_ _02746_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__a31o_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _02062_ _02063_ _02076_ _02081_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__o31a_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08475_ _02014_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__xor2_1
X_07426_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _01143_ VGND
+ VGND VPWR VPWR _01160_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07357_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ _01082_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07288_ _01032_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ _01019_ _01035_ _01026_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09027_ _02312_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] VGND
+ VGND VPWR VPWR _02510_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold250 r_i_alpha1\[12\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold261 _00433_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND VGND VPWR
+ VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03304_ VGND
+ VGND VPWR VPWR _03305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12940_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05915_
+ _05878_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _05862_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__or2_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ clknet_leaf_45_i_clk _00155_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _04957_ _04953_ _04954_ _04754_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__a31o_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11753_ _04895_ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__and2_1
X_14541_ clknet_leaf_38_i_clk _00087_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _03978_ _03988_ _03989_ _03631_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a31o_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__and2b_1
X_14472_ clknet_leaf_7_i_clk _00018_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10635_ _03925_ _03927_ _03928_ _03604_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__a31o_1
X_13423_ _06323_ _06329_ _06327_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13354_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _06269_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10566_ _03861_ _03864_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12305_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05376_ VGND
+ VGND VPWR VPWR _05377_ sky130_fd_sc_hd__xor2_1
X_13285_ _06215_ _06220_ _06201_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10497_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03796_ VGND
+ VGND VPWR VPWR _03805_ sky130_fd_sc_hd__nand2_1
X_15024_ clknet_leaf_97_i_clk _00569_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_12236_ _05142_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05315_
+ _05316_ _05170_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12167_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05254_ VGND
+ VGND VPWR VPWR _05255_ sky130_fd_sc_hd__xnor2_2
X_11118_ _04340_ _04345_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__and2_1
X_12098_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05194_
+ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__and2_1
X_11049_ _04278_ _04280_ _04287_ _04047_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 in_alpha[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14808_ clknet_leaf_67_i_clk _00353_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ clknet_leaf_64_i_clk _00284_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_08260_ _01562_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08191_ _01559_ _01777_ _01453_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07975_ _01576_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__or2b_1
X_09714_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03120_ VGND
+ VGND VPWR VPWR _03121_ sky130_fd_sc_hd__xor2_1
X_09645_ _02748_ _03056_ _03057_ _03058_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _02993_ _02989_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__a21oi_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08527_ _02061_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08458_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[5\] _01992_ _01880_ VGND
+ VGND VPWR VPWR _02003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07409_ _01143_ _01144_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08389_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[14\] _01942_ _01866_
+ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10420_ _03724_ _03727_ _03722_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10351_ _03671_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _03606_
+ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13070_ _05998_ _06035_ _06036_ _05938_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__o211a_1
X_10282_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _03609_
+ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__or2_1
X_12021_ _05130_ net218 _04979_ _05133_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13972_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _06807_ VGND
+ VGND VPWR VPWR _06815_ sky130_fd_sc_hd__or2_1
X_12923_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _05907_
+ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ net645 _05848_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__or2_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _04942_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__or2_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12785_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05781_ VGND
+ VGND VPWR VPWR _05794_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ clknet_leaf_47_i_clk _00070_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.i_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11736_ _04870_ _04877_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__and2_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14455_ clknet_leaf_42_i_clk _00001_ VGND VGND VPWR VPWR r_i_alpha1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _04820_
+ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13406_ _06234_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10618_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03905_ _03650_
+ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__o21a_1
X_11598_ _04756_ net166 _04762_ _04764_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14386_ _07161_ _07155_ _07166_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10549_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03849_ VGND
+ VGND VPWR VPWR _03850_ sky130_fd_sc_hd__xnor2_1
X_13337_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06265_
+ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13268_ _06202_ net295 _06203_ _06208_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__o211a_1
X_15007_ clknet_leaf_103_i_clk _00552_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12219_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05279_ VGND
+ VGND VPWR VPWR _05302_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13199_ _06146_ _06147_ _06150_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_138_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07760_ _01338_ _01406_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__nand2_1
X_07691_ net5 _01355_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__xnor2_1
X_09430_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _02863_ VGND
+ VGND VPWR VPWR _02864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09361_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _02796_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08312_ _01877_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR _01878_ sky130_fd_sc_hd__nand2_1
X_09292_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08243_ _01572_ _01667_ _01820_ _01821_ _01485_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_28_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08174_ _01472_ _01755_ _01762_ _01763_ _01457_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07958_ _01472_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_4
X_07889_ _01329_ _01502_ _01503_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__o21a_1
X_09628_ _03036_ _03029_ _03041_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09559_ _02972_ _02974_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__a21o_1
X_12570_ _05601_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11521_ _04699_ _04695_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11452_ _04442_ _04636_ _04637_ _04456_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__o211a_1
X_14240_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ _07042_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10403_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14171_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06977_
+ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11383_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04565_ _04570_
+ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_150_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13122_ _06071_ _06073_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__or2_1
X_10334_ _03658_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _06010_ _06018_
+ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__a21o_1
X_10265_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__clkbuf_4
X_12004_ _05117_ _05119_ _04757_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__o21a_1
X_10196_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03536_ _03206_
+ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13955_ _06788_ _06789_ _06787_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__a21o_1
X_12906_ _05848_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13886_ _06717_ _06737_ _06739_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__o21a_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05499_ VGND
+ VGND VPWR VPWR _05839_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12768_ _05761_ _05754_ _05774_ _05778_ _05773_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__o32a_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14507_ clknet_leaf_27_i_clk _00053_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_1
X_11719_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04794_ _04864_
+ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12699_ _05707_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _05716_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14438_ _07208_ _07210_ _07213_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__a21oi_1
Xinput10 in_alpha[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
Xinput21 in_x[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 in_x[3] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xinput43 in_y[13] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput54 in_y[7] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14369_ _06911_ net624 _07153_ _07154_ _01456_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__o221a_1
XFILLER_0_110_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08930_ _02412_ _02417_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08861_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _02359_
+ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__or2b_1
X_07812_ net200 _01345_ _01441_ _01442_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a22o_1
X_08792_ _02304_ _02301_ _02305_ _01870_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__o31ai_1
X_07743_ _01393_ _01394_ net239 _01333_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07674_ _00992_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkinv_4
X_09413_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _02850_ sky130_fd_sc_hd__buf_2
XFILLER_0_90_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09344_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02791_
+ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09275_ _02715_ _02728_ _02729_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08226_ _01330_ _01630_ _01529_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08157_ net28 net46 VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08088_ _01664_ _01666_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10050_ _03414_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06607_
+ _06612_ _06584_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__o31ai_1
X_10952_ _04199_ _04200_ _04201_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13671_ _06553_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__buf_2
X_10883_ _04138_ _04139_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__and2_1
X_15410_ clknet_leaf_29_i_clk _00955_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12622_ _05647_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15341_ clknet_leaf_50_i_clk _00886_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_12553_ _05587_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11504_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04684_ VGND
+ VGND VPWR VPWR _04685_ sky130_fd_sc_hd__xnor2_2
X_15272_ clknet_leaf_11_i_clk _00817_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12484_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _05524_ _05529_ _05391_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14223_ _07017_ _07028_ _04961_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11435_ _04237_ _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11366_ _04549_ _04558_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__and2b_1
X_14154_ _06966_ _06969_ _06904_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13105_ _06060_ _06065_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__nor2_1
X_10317_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _03629_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_2_i_clk clknet_4_2_0_i_clk VGND VGND VPWR VPWR clknet_leaf_2_i_clk sky130_fd_sc_hd__clkbuf_16
X_11297_ _04484_ _04491_ _04492_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _06911_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__nand2_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _05848_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _06008_ sky130_fd_sc_hd__or2_1
X_10248_ _03564_ _03579_ _03592_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__and3b_1
XFILLER_0_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10179_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03530_ VGND
+ VGND VPWR VPWR _03531_ sky130_fd_sc_hd__xnor2_2
X_14987_ clknet_leaf_104_i_clk _00532_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_13938_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ _06586_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13869_ _06553_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07390_ _01095_ net230 _01127_ _01128_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09060_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _02525_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08011_ _01609_ _01610_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09962_ _03333_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08913_ _02406_ _02404_ _02405_ _02369_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__a31o_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _03186_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__or2_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02335_
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND VPWR
+ VPWR _02349_ sky130_fd_sc_hd__o21a_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _02277_ _02286_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__nor2_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _00991_ net16 net17 VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__o21a_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07657_ _01330_ _01255_ _01276_ _01331_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_125_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07588_ _01258_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09327_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _02768_
+ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09258_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _02706_ _02704_
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND VPWR VPWR
+ _02719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08209_ _01765_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09189_ _02650_ _02654_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__and2_1
X_11220_ _04378_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11151_ _04378_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__clkbuf_2
X_10102_ _03458_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__nand2_1
X_11082_ _04317_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__nand2_1
X_14910_ clknet_leaf_81_i_clk _00455_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_10033_ _03398_ _03385_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__and2_1
X_14841_ clknet_leaf_85_i_clk _00386_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_14772_ clknet_leaf_52_i_clk _00317_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11984_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05072_ VGND
+ VGND VPWR VPWR _05103_ sky130_fd_sc_hd__and2_1
X_13723_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _06594_
+ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__or2_1
X_10935_ _04184_ _04185_ _03997_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13654_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06514_ VGND
+ VGND VPWR VPWR _06543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10866_ _04113_ _04115_ _04111_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12605_ _05601_ _05633_ _05609_ _05629_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__o211ai_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _06481_ _06482_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__xor2_1
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10797_ _01474_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15324_ clknet_leaf_18_i_clk _00869_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12536_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15255_ clknet_leaf_3_i_clk _00800_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_12467_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05513_
+ _05501_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14206_ _07010_ _07012_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__nand2_1
X_11418_ _04601_ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__xor2_1
X_15186_ clknet_leaf_124_i_clk _00731_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12398_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] net653 _05430_
+ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14137_ _06928_ net334 _06954_ _06955_ _06922_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__o221a_1
X_11349_ _04540_ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14068_ _06893_ _06895_ _06898_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13019_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _05982_ VGND
+ VGND VPWR VPWR _05992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08560_ _02095_ _02096_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__nor2_1
X_07511_ _01010_ _01170_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08491_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\]
+ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__or2_1
X_07442_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07373_ _01095_ net208 _01112_ _01113_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_103_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_103_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09112_ _02580_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _02585_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09043_ _02481_ _02502_ _02519_ _02523_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold410 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold421 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_118_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_118_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold432 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND VGND
+ VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold465 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _00376_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ _03318_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__nor2_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03249_
+ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__or2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _02329_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _02332_ _02334_ _02309_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__o221a_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _02092_ _02274_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__nand2_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _01370_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _02211_ _02212_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__nand2_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ net175 _03999_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__or2_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10651_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03942_ _03651_
+ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10582_ _03862_ _03879_ _03649_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__o21a_1
X_13370_ _06251_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12321_ _05142_ net420 _05389_ _05390_ _05391_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15040_ clknet_leaf_96_i_clk _00585_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_12252_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05291_ VGND
+ VGND VPWR VPWR _05330_ sky130_fd_sc_hd__or2_1
X_11203_ net463 VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__inv_2
X_12183_ _05246_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11134_ _04363_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_82_i_clk clknet_4_7_0_i_clk VGND VGND VPWR VPWR clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11065_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04302_ VGND
+ VGND VPWR VPWR _04303_ sky130_fd_sc_hd__nand2_1
X_10016_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03370_ _03206_
+ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__o21a_1
X_14824_ clknet_leaf_52_i_clk _00369_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_97_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_97_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14755_ clknet_leaf_64_i_clk _00300_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11967_ _05087_ _05088_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13706_ net516 _06582_ _06584_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__o21ai_1
X_10918_ _04153_ _04163_ _04170_ _03994_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_20_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14686_ clknet_leaf_62_i_clk _00231_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11898_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05025_ _04795_
+ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13637_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06514_ VGND
+ VGND VPWR VPWR _06528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10849_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ _04093_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__or3_4
XFILLER_0_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13568_ _06466_ _06467_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15307_ clknet_leaf_23_i_clk _00852_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12519_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05557_
+ _05487_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_35_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13499_ _06405_ _06406_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15238_ clknet_leaf_14_i_clk _00783_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15169_ clknet_leaf_113_i_clk _00714_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07991_ _01577_ _01584_ _01576_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09730_ _03111_ _03135_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09661_ _02634_ _03071_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__nand2_1
X_08612_ _02136_ _02141_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09592_ _03000_ _03009_ _03010_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08543_ _02061_ _02077_ _02079_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08474_ _01998_ _02005_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07425_ _01026_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07356_ _01047_ _01096_ _01097_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07287_ _01033_ _01034_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09026_ _02507_ _02500_ _02503_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold240 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold251 r_i_alpha1\[8\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 diff2\[7\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold273 diff3\[8\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\] VGND VGND VPWR VPWR
+ net401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _03205_ VGND VGND VPWR
+ VPWR _03304_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09859_ _03243_ _03245_ _02850_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__mux2_1
X_12870_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND VPWR
+ VPWR _05863_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _04953_ _04954_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__a21oi_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ clknet_leaf_38_i_clk _00086_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _04894_ VGND
+ VGND VPWR VPWR _04896_ sky130_fd_sc_hd__or2b_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10703_ _03978_ _03988_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__a21oi_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ clknet_leaf_5_i_clk _00017_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _04773_ net391 _04832_ _04833_ _04788_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__o221a_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13422_ _06338_ _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__nand2_1
X_10634_ _03903_ _03910_ _03915_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13353_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _06275_
+ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__or2_1
X_10565_ _03861_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12304_ _05163_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13284_ _06215_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__nor2_1
X_10496_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03796_ _03789_
+ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15023_ clknet_leaf_98_i_clk _00568_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_12235_ _05313_ _05314_ _05129_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a21o_1
X_12166_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05253_ VGND
+ VGND VPWR VPWR _05254_ sky130_fd_sc_hd__xnor2_2
X_11117_ _04348_ _04349_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__and2_1
X_12097_ _04829_ _05191_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__o21a_1
X_11048_ _04278_ _04280_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__a21oi_1
Xinput8 in_alpha[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14807_ clknet_leaf_67_i_clk _00352_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12999_ _05966_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14738_ clknet_leaf_64_i_clk _00283_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14669_ clknet_leaf_54_i_clk _00214_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08190_ _01559_ _01777_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07974_ net50 net32 VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__or2b_1
X_09713_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03107_ _02770_
+ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09644_ _01474_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09575_ _02994_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__and2_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08526_ _02062_ _02063_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08457_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR VPWR
+ _02002_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07408_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _01129_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08388_ _01938_ _01939_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\]
+ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07339_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _01069_ VGND
+ VGND VPWR VPWR _01083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10350_ _03671_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09009_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02492_ VGND
+ VGND VPWR VPWR _02493_ sky130_fd_sc_hd__xor2_2
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10281_ _03607_ net254 _03568_ _03616_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12020_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _05132_
+ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__or2_1
X_13971_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _06807_ VGND
+ VGND VPWR VPWR _06814_ sky130_fd_sc_hd__and2_1
X_12922_ _05567_ _05904_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__o21a_1
X_12853_ _05843_ net204 _05847_ _05850_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__o211a_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04915_ VGND
+ VGND VPWR VPWR _04943_ sky130_fd_sc_hd__and2_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05781_ VGND
+ VGND VPWR VPWR _05793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14523_ clknet_leaf_42_i_clk _00069_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in
+ sky130_fd_sc_hd__dfxtp_1
X_11735_ _04862_ _04879_ _04880_ _04739_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__o211a_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ clknet_leaf_39_i_clk _00000_ VGND VGND VPWR VPWR r_i_alpha1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11666_ _04818_ _04819_ _04795_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13405_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10617_ _03606_ _03911_ _03912_ _03780_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14385_ _06911_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _07167_
+ _07168_ _01456_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__o221a_1
X_11597_ net162 _04758_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13336_ _05928_ _06262_ _06264_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__o21a_1
X_10548_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _03649_ VGND VGND VPWR
+ VPWR _03849_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13267_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] _06205_
+ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__or2_1
X_10479_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03787_ _03788_
+ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15006_ clknet_leaf_103_i_clk _00551_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_12218_ _05301_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
X_13198_ _06148_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__and2_1
X_12149_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _05238_ VGND
+ VGND VPWR VPWR _05239_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07690_ _01355_ _01356_ net181 _01345_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__a2bb2o_1
X_09360_ _02748_ _02803_ _02805_ _02260_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__o211a_1
X_08311_ _01869_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_4
X_09291_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__buf_4
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08242_ _01669_ _01819_ _01472_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08173_ _01748_ _01760_ _01761_ _01329_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07957_ _01539_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\] _01560_ _01561_
+ _01513_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__o221a_1
X_07888_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\] _01498_ _01328_ VGND
+ VGND VPWR VPWR _01503_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09627_ _03036_ _03029_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09558_ _02972_ _02974_ _02967_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08509_ _02049_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _02050_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09489_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11520_ _04695_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11451_ _04444_ net513 VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10402_ _03626_ net393 _03717_ _03718_ _03633_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__o221a_1
X_14170_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06978_
+ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nand2_1
X_11382_ _04431_ net556 _04575_ _04576_ _04539_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13121_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _06080_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10333_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _03644_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__or3_1
X_13052_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _06003_ VGND
+ VGND VPWR VPWR _06021_ sky130_fd_sc_hd__xnor2_1
X_10264_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12003_ _05117_ _05119_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__nand2_1
X_10195_ _03545_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
X_13954_ _06797_ _06798_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__or2b_1
X_12905_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _05892_
+ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__xor2_1
X_13885_ _06721_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12836_ _05836_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__xnor2_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _05759_ _05772_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__nor2_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ clknet_leaf_31_i_clk _00052_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_1
X_11718_ _04794_ _04864_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__a21oi_1
X_12698_ _05713_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14437_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _07156_ VGND
+ VGND VPWR VPWR _07213_ sky130_fd_sc_hd__xor2_1
X_11649_ _04771_ _04805_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__nand2_1
Xinput11 in_alpha[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
Xinput22 in_x[10] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput33 in_x[4] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xinput44 in_y[14] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput55 in_y[8] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
X_14368_ _07146_ _07148_ _07152_ _06926_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__a31o_1
X_13319_ _06204_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14299_ _07092_ _07093_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _06903_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_150_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08860_ _02314_ _02361_ _02362_ _02260_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__o211a_1
X_07811_ _01003_ net7 _01435_ _00993_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__o31a_1
X_08791_ _02304_ _02301_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__o21a_1
X_07742_ net4 _01391_ _01344_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__a21oi_1
X_07673_ _01343_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
X_09412_ _02844_ net474 _02848_ _02849_ _02827_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__o221a_1
X_09343_ _02789_ _02790_ _02772_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09274_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _02726_ VGND
+ VGND VPWR VPWR _02733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08225_ _01805_ _01806_ _01562_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08156_ net46 net28 VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08087_ net22 net40 VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08989_ _02473_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10951_ _03997_ net554 _01794_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13670_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__buf_2
X_10882_ _04128_ _04129_ _04131_ _04137_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__a31o_1
X_12621_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _05648_ _05643_
+ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15340_ clknet_leaf_50_i_clk _00885_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12552_ _05290_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11503_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04683_ VGND
+ VGND VPWR VPWR _04684_ sky130_fd_sc_hd__xor2_2
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15271_ clknet_leaf_12_i_clk _00816_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12483_ _05526_ _05527_ _05528_ _05490_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__o31ai_1
X_14222_ _07025_ _07026_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11434_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04620_ VGND
+ VGND VPWR VPWR _04621_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14153_ _06967_ _06968_ _06934_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11365_ _04431_ _04557_ _04560_ _04561_ _04539_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13104_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _06064_ VGND
+ VGND VPWR VPWR _06065_ sky130_fd_sc_hd__xnor2_1
X_10316_ _03625_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _03641_ _03643_ _03633_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14084_ _06909_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__clkbuf_4
X_11296_ _04478_ _04479_ _04497_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__o21a_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _06005_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__nor2_1
X_10247_ _03583_ _03588_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__nor2_1
X_10178_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03529_ VGND
+ VGND VPWR VPWR _03530_ sky130_fd_sc_hd__xor2_2
X_14986_ clknet_leaf_104_i_clk _00531_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_13937_ _06555_ _06782_ _06783_ _06747_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13868_ _06721_ _06722_ _06723_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12819_ _05486_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05822_
+ _05823_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13799_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _06661_ VGND
+ VGND VPWR VPWR _06663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08010_ net35 _01608_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09961_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03332_ VGND
+ VGND VPWR VPWR _03334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08912_ _02404_ _02405_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _03271_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__xnor2_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _02330_
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND VPWR
+ VPWR _02348_ sky130_fd_sc_hd__a21o_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08774_ _01924_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] VGND
+ VGND VPWR VPWR _02290_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07725_ net196 _01333_ _01380_ _01381_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__o22a_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07656_ net178 _01255_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07587_ diff2\[4\] _01270_ _01272_ diff3\[4\] _01274_ VGND VGND VPWR VPWR _01275_
+ sky130_fd_sc_hd__a221o_1
X_09326_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND VPWR
+ VPWR _02776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09257_ _02698_ _02705_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08208_ _01572_ _01592_ _01791_ _01792_ _01457_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09188_ _02650_ _02654_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08139_ _01703_ _01728_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__a21boi_1
X_11150_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _04378_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10101_ _03446_ _03451_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__a21o_1
X_11081_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04316_ VGND
+ VGND VPWR VPWR _04318_ sky130_fd_sc_hd__or2_1
X_10032_ _03398_ _03385_ _03383_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__o21a_1
X_14840_ clknet_leaf_84_i_clk _00385_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14771_ clknet_leaf_52_i_clk _00316_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11983_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05072_ VGND
+ VGND VPWR VPWR _05102_ sky130_fd_sc_hd__nor2_1
X_13722_ _06561_ net490 _06485_ _06598_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__o211a_1
X_10934_ _04184_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13653_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06514_ VGND
+ VGND VPWR VPWR _06542_ sky130_fd_sc_hd__or2_1
X_10865_ _04121_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__nand2_1
X_12604_ _05608_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _06472_ _06475_ _06471_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__o21a_1
X_10796_ _03999_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ clknet_leaf_18_i_clk _00868_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12535_ _05521_ net471 _05570_ _05571_ _05544_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__o221a_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15254_ clknet_leaf_5_i_clk _00799_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_12466_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05513_
+ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14205_ _06999_ _07003_ _07011_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__o21ai_2
X_11417_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _04605_ VGND
+ VGND VPWR VPWR _04606_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15185_ clknet_leaf_123_i_clk _00730_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12397_ _05142_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05458_
+ _05459_ _05391_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_13_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_14136_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06953_
+ _01862_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__o21ai_1
X_11348_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04541_ _04545_
+ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14067_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06845_ VGND
+ VGND VPWR VPWR _06898_ sky130_fd_sc_hd__xor2_1
X_11279_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04482_ VGND
+ VGND VPWR VPWR _04483_ sky130_fd_sc_hd__xor2_1
X_13018_ _05991_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14969_ clknet_leaf_105_i_clk _00514_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_07510_ _01016_ net229 _01225_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08490_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _02031_
+ _02032_ _01908_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07441_ _01019_ _01170_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07372_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09111_ _02329_ net325 _02381_ _02584_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09042_ _02520_ _02515_ _02521_ _02500_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_143_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold400 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND VPWR VPWR
+ net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold433 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND VGND VPWR
+ VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold477 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND VGND VPWR
+ VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _03317_ VGND
+ VGND VPWR VPWR _03319_ sky130_fd_sc_hd__nor2_1
Xhold488 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND VGND
+ VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND VGND VPWR
+ VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _02850_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__nand2_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _02327_ _02330_ _02331_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__a31o_1
X_08757_ _02092_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__or2_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ net362 _01369_ _01358_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__mux2_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _02025_ _02210_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__nand2_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ diff2\[14\] _01269_ _01271_ diff3\[14\] _01316_ VGND VGND VPWR VPWR _01317_
+ sky130_fd_sc_hd__a221o_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_i_clk clknet_4_0_0_i_clk VGND VGND VPWR VPWR clknet_leaf_1_i_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10650_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03941_ VGND
+ VGND VPWR VPWR _03942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09309_ _02409_ _02758_ _02759_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10581_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12320_ _04538_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12251_ _05142_ net594 _05328_ _05329_ _05170_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__o221a_1
X_11202_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _04398_ _04414_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a31o_1
X_12182_ _05234_ _05267_ _05268_ _05080_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__o211a_1
X_11133_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04338_ VGND
+ VGND VPWR VPWR _04364_ sky130_fd_sc_hd__nand2_1
X_11064_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04301_ VGND
+ VGND VPWR VPWR _04302_ sky130_fd_sc_hd__xnor2_1
X_10015_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03372_ VGND
+ VGND VPWR VPWR _03383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14823_ clknet_leaf_16_i_clk _00368_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11966_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05081_ _05085_
+ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14754_ clknet_leaf_64_i_clk _00299_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10917_ _04153_ _04163_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__a21oi_1
X_13705_ _06562_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__clkbuf_4
X_14685_ clknet_leaf_62_i_clk _00230_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11897_ _04557_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND VGND VPWR VPWR
+ _05025_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13636_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06488_ VGND
+ VGND VPWR VPWR _06527_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10848_ _04048_ _04106_ _04107_ _04063_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13567_ _06450_ _06456_ _06454_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__o21ba_1
X_10779_ _03993_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12518_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05557_
+ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15306_ clknet_leaf_23_i_clk _00851_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13498_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06351_ VGND
+ VGND VPWR VPWR _06406_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12449_ _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__clkbuf_4
X_15237_ clknet_leaf_12_i_clk _00782_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15168_ clknet_leaf_113_i_clk net351 VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14119_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _06917_ VGND VGND
+ VPWR VPWR _06940_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15099_ clknet_leaf_118_i_clk _00644_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_07990_ _01589_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09660_ _02634_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__or2_1
X_08611_ _02136_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__nor2_1
X_09591_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _02986_ VGND
+ VGND VPWR VPWR _03010_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08542_ _02078_ _02072_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08473_ _02015_ _02004_ _02016_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07424_ _01044_ net177 _01158_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07355_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _01077_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07286_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] VGND VGND VPWR VPWR
+ _01034_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09025_ _02500_ _02503_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold230 diff1\[6\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND
+ VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 net93 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 diff1\[2\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _00142_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _01248_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _03303_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_1
X_09858_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__inv_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _02319_ sky130_fd_sc_hd__clkbuf_4
X_09789_ _03184_ net145 _03017_ _03187_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__o211a_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _04955_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__or2_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _04894_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _04895_ sky130_fd_sc_hd__or2b_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _03944_ VGND
+ VGND VPWR VPWR _03989_ sky130_fd_sc_hd__xor2_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ clknet_leaf_5_i_clk _00016_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11682_ _04831_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _04755_
+ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _06333_ _06337_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__a21o_1
X_10633_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03914_ _03926_
+ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_107_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13352_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _06277_ _06278_ _06197_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__o221a_1
XFILLER_0_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10564_ _03752_ _03863_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12303_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__or4_2
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13283_ _06218_ _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10495_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03796_ _03792_
+ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__o21ai_1
X_15022_ clknet_leaf_97_i_clk _00567_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12234_ _05313_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nor2_1
X_12165_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ net121 _05163_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__o31a_1
XFILLER_0_102_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11116_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04338_ VGND
+ VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nand2_1
X_12096_ _04829_ _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11047_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_102_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_102_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput9 in_alpha[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
XFILLER_0_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14806_ clknet_leaf_66_i_clk _00351_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_12998_ _05971_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_117_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_117_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14737_ clknet_leaf_64_i_clk _00282_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_11949_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _05069_ VGND
+ VGND VPWR VPWR _05073_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ clknet_leaf_54_i_clk _00213_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13619_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _06511_
+ _06512_ _06285_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14599_ clknet_leaf_44_i_clk _00144_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07973_ net32 net50 VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__and2b_1
X_09712_ _03119_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
X_09643_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _03057_ sky130_fd_sc_hd__or2_1
X_09574_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _02986_ VGND
+ VGND VPWR VPWR _02995_ sky130_fd_sc_hd__or2_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _02037_ _02064_ _02051_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08456_ _01998_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_81_i_clk clknet_4_6_0_i_clk VGND VGND VPWR VPWR clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07407_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ _01129_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__or3_4
XFILLER_0_46_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08387_ _01891_ net628 _01940_ _01941_ _01908_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07338_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _01069_ VGND
+ VGND VPWR VPWR _01082_ sky130_fd_sc_hd__or2_4
XFILLER_0_104_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07269_ _01017_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09008_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _02483_ _02343_
+ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10280_ net234 _03609_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13970_ _06555_ _06812_ _06813_ _06747_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__o211a_1
X_12921_ _05567_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_34_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ net646 _05848_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__or2_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04930_ VGND
+ VGND VPWR VPWR _04942_ sky130_fd_sc_hd__nor2_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _05632_ _05791_ _05792_ _05675_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__o211a_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11734_ _04765_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _04880_ sky130_fd_sc_hd__or2_1
X_14522_ clknet_leaf_2_i_clk _00068_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11665_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04807_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14453_ _07059_ _07225_ _07226_ _01475_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10616_ _03608_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _03912_ sky130_fd_sc_hd__or2_1
X_13404_ _06317_ _06319_ _06316_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14384_ _07160_ _07162_ _07166_ _06926_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__a31o_1
X_11596_ _04756_ net151 _04762_ _04763_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13335_ _05928_ _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10547_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _03848_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13266_ _06202_ net140 _06203_ _06207_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__o211a_1
X_10478_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03773_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__or3b_1
X_15005_ clknet_leaf_103_i_clk net464 VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12217_ _05290_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13197_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06136_ VGND
+ VGND VPWR VPWR _06149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12148_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05237_ VGND
+ VGND VPWR VPWR _05238_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12079_ _04829_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _05171_ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08310_ _01869_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_4
X_09290_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08241_ _01669_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08172_ _01760_ _01761_ _01748_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput110 net110 VGND VGND VPWR VPWR out_sintheta[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07956_ net21 _01472_ _01559_ _01453_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__a31o_1
X_07887_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] _01487_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[7\] VGND VGND VPWR VPWR _01502_
+ sky130_fd_sc_hd__o211a_1
X_09626_ _03039_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09557_ _02844_ net636 _02978_ _02979_ _02827_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08508_ _02047_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09488_ _02844_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _02915_
+ _02916_ _02827_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08439_ _01984_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11450_ _04631_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10401_ _03714_ _03716_ _03642_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11381_ _04568_ _04570_ _04574_ _04396_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13120_ _06079_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
X_10332_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03634_ VGND VGND
+ VPWR VPWR _03657_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13051_ _06014_ _06020_ _04961_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10263_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__clkbuf_4
X_12002_ _04903_ _05081_ _05092_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__a22o_1
X_10194_ _03535_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13953_ _06794_ _06796_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__nand2_1
X_12904_ _05567_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _05884_ _05891_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__a31o_1
X_13884_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _06716_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__o21a_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05789_ VGND
+ VGND VPWR VPWR _05837_ sky130_fd_sc_hd__xnor2_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _05500_ net264 _05495_ _05777_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14505_ clknet_leaf_27_i_clk _00051_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_1
X_11717_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__or4_2
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _05359_ _05712_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11648_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _04804_
+ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__xnor2_1
X_14436_ _07203_ _07212_ _01766_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_126_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 in_alpha[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 in_x[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput34 in_x[5] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput45 in_y[15] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
XFILLER_0_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11579_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04378_ VGND
+ VGND VPWR VPWR _04752_ sky130_fd_sc_hd__or2_1
X_14367_ _07146_ _07148_ _07152_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__a21oi_1
Xinput56 in_y[9] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13318_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _06249_
+ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14298_ _07089_ _07091_ _07088_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13249_ _05978_ _06142_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07810_ _01003_ _01435_ net7 VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__o21ai_2
X_08790_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[17\] _02298_ VGND VGND VPWR
+ VPWR _02305_ sky130_fd_sc_hd__xnor2_1
X_07741_ net4 _01391_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07672_ net347 _01342_ _01000_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__mux2_1
X_09411_ _02847_ _02845_ _02846_ _02761_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09342_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _02777_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09273_ _02322_ net579 _02731_ _02732_ _02689_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08224_ _01609_ _01627_ _01801_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08155_ _01717_ net446 _01635_ _01745_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08086_ _01679_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__nor2_2
XFILLER_0_113_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08988_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _02471_ VGND
+ VGND VPWR VPWR _02474_ sky130_fd_sc_hd__and2b_1
X_07939_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[16\] _01545_ _01480_
+ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10950_ _04189_ _04194_ _04198_ _03997_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09609_ _03019_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _03025_ sky130_fd_sc_hd__and2b_1
X_10881_ _04128_ _04129_ _04131_ _04137_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__nand4_1
X_12620_ _05641_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12551_ _05584_ _05585_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ _05486_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11502_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04671_ _04413_
+ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__o21a_1
X_12482_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05507_ VGND VGND
+ VPWR VPWR _05528_ sky130_fd_sc_hd__and4_1
X_15270_ clknet_leaf_11_i_clk _00815_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11433_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _04412_ VGND VGND VPWR
+ VPWR _04620_ sky130_fd_sc_hd__o31a_1
X_14221_ _07025_ _07026_ _01862_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14152_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06960_
+ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11364_ _04558_ _04559_ _04391_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13103_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06063_ VGND
+ VGND VPWR VPWR _06064_ sky130_fd_sc_hd__xnor2_1
X_10315_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03640_
+ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14083_ _06909_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__buf_4
X_11295_ _04486_ _04493_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__nor2_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _06004_ _06000_ _06002_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__and3_1
X_10246_ _03201_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] VGND
+ VGND VPWR VPWR _03591_ sky130_fd_sc_hd__and2_1
X_10177_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03521_ _03206_
+ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14985_ clknet_leaf_105_i_clk _00530_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_13936_ _06732_ net578 VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13867_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _06707_ VGND
+ VGND VPWR VPWR _06723_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12818_ _05821_ _05816_ _05818_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__o31a_1
X_13798_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _06661_ VGND
+ VGND VPWR VPWR _06662_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _05753_ _05754_ _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__a21o_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14419_ _06909_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _07198_ sky130_fd_sc_hd__or2_1
X_15399_ clknet_leaf_30_i_clk _00944_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09960_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03332_ VGND
+ VGND VPWR VPWR _03333_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08911_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR _02406_ sky130_fd_sc_hd__inv_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09891_ _03207_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _03267_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__o211a_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _02329_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _02346_ _02347_ _02309_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__o221a_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _01877_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _02288_
+ _02289_ _02055_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07724_ _00991_ net16 _00993_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__o21ai_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07586_ _01273_ diff1\[4\] VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09325_ _02757_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _02774_ _02775_ _02689_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09256_ _02715_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08207_ _01589_ _01790_ _01470_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09187_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02653_ VGND
+ VGND VPWR VPWR _02654_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08138_ _01690_ _01729_ _01706_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ net38 net56 VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__and2_1
X_10100_ _03450_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _03459_ sky130_fd_sc_hd__and2b_1
X_11080_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04316_ VGND
+ VGND VPWR VPWR _04317_ sky130_fd_sc_hd__nand2_1
X_10031_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR
+ VPWR _03398_ sky130_fd_sc_hd__inv_2
X_14770_ clknet_leaf_52_i_clk _00315_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11982_ _04862_ _05100_ _05101_ _05080_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13721_ _06563_ _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__nand2_1
X_10933_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04177_ _04179_
+ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10864_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _04120_ VGND
+ VGND VPWR VPWR _04122_ sky130_fd_sc_hd__or2b_1
X_13652_ _06324_ _06514_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12603_ _05487_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__buf_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10795_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _04061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _06479_ _06480_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15322_ clknet_leaf_18_i_clk _00867_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _05569_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _05487_
+ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__a21o_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15253_ clknet_leaf_3_i_clk _00798_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_12465_ _05203_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _05504_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14204_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _07002_ VGND
+ VGND VPWR VPWR _07011_ sky130_fd_sc_hd__nand2_1
X_11416_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04604_ VGND
+ VGND VPWR VPWR _04605_ sky130_fd_sc_hd__xnor2_1
X_15184_ clknet_leaf_124_i_clk _00729_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12396_ _05456_ _05457_ _05129_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11347_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14135_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06953_
+ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11278_ _04413_ _04481_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__nand2_1
X_14066_ _06888_ _06897_ _04961_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__o21a_1
X_13017_ _05990_ _01512_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__and2b_1
X_10229_ _03561_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__nand2_1
X_14968_ clknet_leaf_95_i_clk _00513_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13919_ _06501_ _06768_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__and2_1
X_14899_ clknet_leaf_87_i_clk _00444_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_07440_ _01171_ _01022_ _01023_ _01172_ _01026_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07371_ _01076_ _01107_ _01111_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09110_ _02582_ _02583_ _02320_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09041_ _02520_ _02515_ _02513_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold401 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND VGND
+ VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold412 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold423 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold434 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[14\] VGND VGND VPWR VPWR
+ net551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold456 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold489 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _03317_ VGND
+ VGND VPWR VPWR _03318_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _03237_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _03256_ _03257_ _03258_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__o221a_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _02312_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__buf_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\] _02273_ VGND VGND VPWR
+ VPWR _02274_ sky130_fd_sc_hd__xnor2_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07707_ net9 _01366_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__xnor2_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _02025_ _02210_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ diff2\[17\] diff1\[14\] VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07569_ diff2\[17\] diff1\[17\] VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09308_ _02746_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__buf_4
X_10580_ _03877_ _03874_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09239_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _02702_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12250_ _05326_ _05327_ _05129_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11201_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04407_
+ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__o21ai_1
X_12181_ _05132_ net517 VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__or2_1
X_11132_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04338_ VGND
+ VGND VPWR VPWR _04363_ sky130_fd_sc_hd__or2_1
X_11063_ _03801_ _04192_ net115 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a31o_1
X_10014_ _03382_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__clkbuf_1
X_14822_ clknet_leaf_16_i_clk _00367_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_14753_ clknet_leaf_64_i_clk _00298_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_11965_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05081_ VGND
+ VGND VPWR VPWR _05087_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13704_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _06582_
+ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__and2_1
X_10916_ _04168_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14684_ clknet_leaf_62_i_clk _00229_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_11896_ _04862_ _05023_ _05024_ _04739_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13635_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06524_
+ _06525_ _06526_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__o221a_1
X_10847_ _04010_ net543 VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13566_ _06464_ _06465_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10778_ _04011_ net538 _04003_ _04046_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__o211a_1
X_15305_ clknet_leaf_9_i_clk _00850_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12517_ _05555_ _05556_ _05526_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13497_ _06396_ _06400_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15236_ clknet_leaf_14_i_clk _00781_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12448_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05499_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15167_ clknet_leaf_111_i_clk _00712_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12379_ _05444_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14118_ _06928_ net339 _06938_ _06939_ _06922_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__o221a_1
X_15098_ clknet_leaf_118_i_clk _00643_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_157_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14049_ _06882_ _01512_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08610_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\] _02140_ VGND VGND VPWR
+ VPWR _02141_ sky130_fd_sc_hd__xnor2_1
X_09590_ _03001_ _03005_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__or2b_1
X_08541_ _02078_ _02072_ _02059_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08472_ _02015_ _02004_ _01995_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07423_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _01045_ _01153_
+ _01157_ _01059_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07354_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ _01077_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07285_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR VPWR
+ _01033_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09024_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02506_ VGND
+ VGND VPWR VPWR _02507_ sky130_fd_sc_hd__xor2_2
XFILLER_0_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold220 diff1\[11\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 net104 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 net75 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 diff1\[16\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold286 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR
+ VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _03302_ _03118_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__and2b_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _03238_
+ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__or2_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _02314_ net147 _01945_ _02318_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__o211a_1
X_09788_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _03186_
+ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__or2_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _01869_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _02259_ sky130_fd_sc_hd__or2_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04893_ VGND
+ VGND VPWR VPWR _04894_ sky130_fd_sc_hd__xor2_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _03979_ _03984_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__or2_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _04831_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _04832_ sky130_fd_sc_hd__nor2_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _06333_ _06337_
+ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__nand3_2
XFILLER_0_107_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10632_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03907_ _03914_
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND VGND VPWR VPWR
+ _03926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10563_ _03650_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__nand2_1
X_13351_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _06276_
+ _06216_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12302_ _05366_ _05370_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10494_ _03642_ _03801_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__nor2_1
X_13282_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND VPWR
+ VPWR _06219_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15021_ clknet_leaf_98_i_clk _00566_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12233_ _05307_ _05310_ _05306_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12164_ _05247_ _05249_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11115_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04338_ VGND
+ VGND VPWR VPWR _04348_ sky130_fd_sc_hd__or2_1
X_12095_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05182_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__and3_1
X_11046_ _04284_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__or2b_1
X_14805_ clknet_leaf_67_i_clk _00350_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12997_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _05970_ VGND
+ VGND VPWR VPWR _05972_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14736_ clknet_leaf_65_i_clk _00281_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11948_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14667_ clknet_leaf_54_i_clk _00212_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11879_ _05001_ _04994_ _05007_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13618_ _06503_ _06509_ _06510_ _06200_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14598_ clknet_leaf_44_i_clk _00143_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13549_ _06444_ _06446_ _06443_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15219_ clknet_leaf_15_i_clk _00764_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_i_clk clknet_4_0_0_i_clk VGND VGND VPWR VPWR clknet_leaf_0_i_clk sky130_fd_sc_hd__clkbuf_16
X_07972_ _01463_ net459 _01460_ _01575_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__o211a_1
X_09711_ _03117_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__and2b_1
X_09642_ _03054_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__nor2_1
X_09573_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _02986_ VGND
+ VGND VPWR VPWR _02994_ sky130_fd_sc_hd__nand2_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _02049_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _02064_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08455_ _01876_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _01945_
+ _02000_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07406_ _01044_ net170 _01142_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08386_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\] _01938_ _01939_
+ _01924_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07337_ _01037_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07268_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR _01017_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09007_ _02321_ net616 _02381_ _02491_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09909_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03286_ VGND
+ VGND VPWR VPWR _03287_ sky130_fd_sc_hd__xnor2_1
X_12920_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _05895_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _05843_ net207 _05847_ _05849_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__o211a_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _04935_ _04937_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__and3_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _05792_ sky130_fd_sc_hd__or2_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ clknet_leaf_32_i_clk _00067_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _04877_ _04878_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__xnor2_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06909_ VGND
+ VGND VPWR VPWR _07226_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11664_ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13403_ _06322_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
X_10615_ _03903_ _03910_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14383_ _07160_ _07162_ _07166_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a21oi_1
X_11595_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] _04758_
+ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13334_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _06253_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__and3_1
X_10546_ _03847_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ net648 _06205_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__or2_1
X_10477_ _03786_ _03651_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15004_ clknet_leaf_103_i_clk net461 VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12216_ _05298_ _05299_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _05128_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13196_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06136_ VGND
+ VGND VPWR VPWR _06148_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12147_ _05163_ net121 VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12078_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05177_
+ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__nor2_1
X_11029_ _03669_ net115 VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14719_ clknet_leaf_53_i_clk _00264_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08240_ _01673_ _01810_ _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08171_ _01720_ _01736_ _01735_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput100 net100 VGND VGND VPWR VPWR out_sintheta[15] sky130_fd_sc_hd__clkbuf_4
Xoutput111 net111 VGND VGND VPWR VPWR out_sintheta[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07955_ net21 _01556_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__a21oi_1
X_07886_ _01467_ net629 _01500_ _01501_ _01475_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__o221a_1
X_09625_ _02595_ _03038_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__and2_1
X_09556_ _02975_ _02977_ _02747_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08507_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\] _02034_ _01880_ VGND
+ VGND VPWR VPWR _02048_ sky130_fd_sc_hd__o21a_1
X_09487_ _02905_ _02908_ _02914_ _02761_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08438_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\] _01983_ VGND VGND VPWR
+ VPWR _01985_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08369_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND VPWR
+ VPWR _01926_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_101_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10400_ _03714_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__and2_1
X_11380_ _04568_ _04570_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10331_ _03625_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _03655_ _03656_ _03633_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13050_ _06018_ _06019_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__nor2_1
X_10262_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _03604_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_116_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_116_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12001_ _05104_ _05105_ _05112_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__and3_1
X_10193_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _03543_ _03185_
+ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13952_ _06794_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12903_ _05566_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__nor2_1
X_13883_ _06715_ _06723_ _06729_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__or3_1
X_12834_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05789_ _05829_
+ _05832_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__a22o_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _05774_ _05775_ _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ clknet_leaf_27_i_clk _00050_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
X_11716_ _04853_ _04856_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__or2_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12696_ _05359_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14435_ _07210_ _07211_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__nand2_1
X_11647_ _04801_ _04803_ _04795_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 in_alpha[2] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_126_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput24 in_x[12] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
X_14366_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _07144_ VGND
+ VGND VPWR VPWR _07152_ sky130_fd_sc_hd__xor2_1
XFILLER_0_141_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput35 in_x[6] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput46 in_y[16] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
X_11578_ _04749_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13317_ _05928_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _06241_ _06248_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__a31o_1
X_10529_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03831_ VGND
+ VGND VPWR VPWR _03832_ sky130_fd_sc_hd__xnor2_1
X_14297_ _07088_ _07089_ _07091_ _01861_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__o31ai_1
X_13248_ _06186_ _06189_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13179_ _06117_ _06130_ _06131_ _06132_ _06125_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__a32oi_4
X_07740_ net195 _01338_ _01390_ _01392_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07671_ _01334_ _01341_ _01339_ net17 VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09410_ _02845_ _02846_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_95_i_clk clknet_4_5_0_i_clk VGND VGND VPWR VPWR clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09341_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09272_ _02715_ _02723_ _02728_ _02729_ _02313_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__a41o_1
XFILLER_0_74_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08223_ _01609_ _01801_ _01627_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08154_ _01556_ _01740_ _01744_ _01454_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08085_ net23 net41 VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_i_clk clknet_4_9_0_i_clk VGND VGND VPWR VPWR clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08987_ _02472_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__inv_2
X_07938_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[16\] _01545_ VGND VGND
+ VPWR VPWR _01546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07869_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[5\] _01476_ VGND VGND
+ VPWR VPWR _01487_ sky130_fd_sc_hd__and2_1
X_09608_ _01765_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__clkbuf_4
X_10880_ _04135_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09539_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12550_ _05581_ _05583_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11501_ _04442_ _04681_ _04682_ _04456_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12481_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _05507_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR _05527_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_65_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14220_ _07010_ _07012_ _07009_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11432_ _04619_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__clkbuf_1
X_14151_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06961_
+ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__and2_1
X_11363_ _04558_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__and2_1
X_13102_ _05566_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND
+ VGND VPWR VPWR _06063_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10314_ _03608_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14082_ _01861_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__buf_2
X_11294_ _04442_ _04495_ _04496_ _04456_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__o211a_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _06000_ _06002_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__a21oi_2
X_10245_ _03183_ _03589_ _03590_ _03515_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10176_ _03389_ _03527_ _03528_ _03515_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__o211a_1
X_14984_ clknet_leaf_104_i_clk _00529_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13935_ _06774_ _06781_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__xor2_1
X_13866_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _06716_ _06717_
+ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12817_ _05816_ _05818_ _05821_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13797_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06660_ VGND
+ VGND VPWR VPWR _06661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12748_ _05759_ _05760_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__or2_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12679_ _05699_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14418_ _07193_ _07196_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15398_ clknet_leaf_31_i_clk _00943_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14349_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _07136_ VGND
+ VGND VPWR VPWR _07137_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08910_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _02393_ _02344_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__a31o_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _03264_ _03265_ _02850_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__a21o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _02340_
+ _02345_ _02333_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__a31o_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _02286_ _02287_ _01924_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__a21o_1
X_07723_ _00991_ net16 VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__and2_1
X_07654_ _01328_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07585_ diff2\[17\] VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09324_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _02773_
+ _02747_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09255_ _02711_ _02714_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08206_ _01589_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__nor2_1
X_09186_ _02342_ _02652_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08137_ net25 net43 VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08068_ _01662_ _01663_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10030_ _03373_ _03386_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__nand2_1
X_11981_ _04770_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND
+ VGND VPWR VPWR _05101_ sky130_fd_sc_hd__or2_1
X_13720_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _06596_
+ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__xnor2_1
X_10932_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04177_ VGND
+ VGND VPWR VPWR _04184_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13651_ _06492_ _06517_ _06539_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__nand3_1
X_10863_ _04120_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _04121_ sky130_fd_sc_hd__or2b_1
X_12602_ _05521_ net399 _05630_ _05631_ _05544_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _06463_ VGND
+ VGND VPWR VPWR _06480_ sky130_fd_sc_hd__nand2_1
X_10794_ net651 _04055_ _04054_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__a21oi_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ clknet_leaf_22_i_clk _00866_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12533_ _05569_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _05570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15252_ clknet_leaf_5_i_clk _00797_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_12464_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05507_
+ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _07008_ _07009_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15183_ clknet_leaf_115_i_clk _00728_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12395_ _05456_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14134_ _06647_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _06946_ _06952_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__o31a_1
X_11346_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04543_ _04413_
+ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14065_ _06557_ _06895_ _06896_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__and3_1
X_11277_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__or4_2
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13016_ _05841_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05988_
+ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__o2bb2a_1
X_10228_ _03572_ _03573_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10159_ _03511_ _03512_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__xor2_1
X_14967_ clknet_leaf_95_i_clk _00512_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13918_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06767_ _06553_
+ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__mux2_1
X_14898_ clknet_leaf_87_i_clk _00443_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13849_ _06684_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07370_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _01080_ _01081_
+ _01110_ _01085_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09040_ _02507_ _02516_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_7_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_7_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold413 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold424 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND VGND
+ VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09942_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03316_ VGND
+ VGND VPWR VPWR _03317_ sky130_fd_sc_hd__xor2_1
Xhold479 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR VPWR
+ net596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _02308_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__clkbuf_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _02330_ _02331_ _02327_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__a21oi_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\]
+ _02249_ _01881_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__o31a_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _01366_ _01368_ net188 _01345_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08686_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\] _02209_ VGND VGND VPWR
+ VPWR _02210_ sky130_fd_sc_hd__xor2_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _01315_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ _01261_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09307_ _02758_ _02759_ _02409_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a21oi_2
X_07499_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _01081_ _01057_
+ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09238_ _02699_ _02700_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09169_ _02637_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11200_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12180_ _05265_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__xnor2_1
X_11131_ _04149_ _04338_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11062_ _04011_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _04219_
+ _04300_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__o211a_1
X_10013_ _03024_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__and2_1
X_14821_ clknet_leaf_16_i_clk _00366_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14752_ clknet_leaf_64_i_clk _00297_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11964_ _04769_ net545 _04979_ _05086_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13703_ _06580_ _06581_ _06292_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__mux2_1
X_10915_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04166_ _04167_
+ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__nand3_1
XFILLER_0_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14683_ clknet_leaf_63_i_clk _00228_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_11895_ _04765_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _05024_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13634_ _01474_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__clkbuf_4
X_10846_ _04104_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__xor2_1
X_13565_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _06461_ _06463_
+ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10777_ _04012_ _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15304_ clknet_leaf_22_i_clk _00849_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12516_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05549_
+ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13496_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06352_ VGND
+ VGND VPWR VPWR _06404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15235_ clknet_leaf_11_i_clk _00780_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12447_ _05488_ net169 _05495_ _05498_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15166_ clknet_leaf_110_i_clk _00711_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12378_ _05290_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14117_ _06937_ _06935_ _06936_ _06926_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__a31o_1
X_11329_ _04526_ _04527_ _04523_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15097_ clknet_leaf_117_i_clk _00642_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14048_ _06875_ _06881_ _06562_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__mux2_1
X_08540_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR VPWR
+ _02078_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08471_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR VPWR
+ _02015_ sky130_fd_sc_hd__inv_2
X_07422_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _01051_ _01052_
+ _01156_ _01057_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07353_ _01015_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07284_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _01032_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09023_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _02505_ VGND
+ VGND VPWR VPWR _02506_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold210 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold221 r_i_alpha1\[11\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold232 _01238_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold243 diff1\[1\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 net58 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold265 diff3\[11\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 diff1\[3\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _03201_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _03300_
+ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__a22oi_1
Xhold298 net63 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _03228_ VGND VGND
+ VPWR VPWR _03243_ sky130_fd_sc_hd__and4_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__or2_1
X_09787_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__clkbuf_4
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _02252_ _02257_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__xnor2_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _02189_ _02190_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__o21ai_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _03987_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR _04831_ sky130_fd_sc_hd__inv_2
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10631_ _03923_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13350_ net568 _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10562_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__or4_4
XFILLER_0_134_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12301_ _05373_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13281_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND VPWR
+ VPWR _06218_ sky130_fd_sc_hd__and3_1
X_10493_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] VGND VGND VPWR
+ VPWR _03801_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15020_ clknet_leaf_92_i_clk _00565_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_12232_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05279_ VGND
+ VGND VPWR VPWR _05313_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12163_ _05153_ net484 _05250_ _05251_ _05170_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11114_ _04012_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04346_
+ _04347_ _04059_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__o221a_1
X_12094_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05177_ VGND VGND
+ VPWR VPWR _05191_ sky130_fd_sc_hd__or4_1
X_11045_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04283_ VGND
+ VGND VPWR VPWR _04285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14804_ clknet_leaf_74_i_clk _00349_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12996_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _05970_ VGND
+ VGND VPWR VPWR _05971_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11947_ _05070_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR VPWR
+ _05071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14735_ clknet_leaf_62_i_clk _00280_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14666_ clknet_leaf_54_i_clk _00211_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11878_ _05001_ _04994_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13617_ _06503_ _06509_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10829_ _03976_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14597_ clknet_leaf_44_i_clk net402 VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13548_ _06449_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13479_ _06383_ _06388_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15218_ clknet_leaf_114_i_clk _00763_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15149_ clknet_leaf_125_i_clk _00694_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07971_ _01562_ _01568_ _01574_ _01485_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__o211ai_2
X_09710_ _01765_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09641_ _03039_ _03043_ _03053_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__nor3_1
XFILLER_0_117_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09572_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02987_ VGND
+ VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08523_ _02039_ _02052_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08454_ _01998_ _01999_ _01877_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__o21ai_1
X_07405_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _01045_ _01139_
+ _01141_ _01059_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08385_ _01938_ _01939_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\]
+ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07336_ _01017_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07267_ _01015_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_4
X_09006_ _02489_ _02490_ _02333_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09908_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__and2b_1
X_09839_ _03207_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__nand2_1
X_12850_ net140 _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__or2_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04901_ _04902_ _04938_ _04939_ _04909_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__o2111ai_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05788_ _05790_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__xnor2_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ clknet_leaf_33_i_clk _00066_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11732_ _04863_ _04870_ _04868_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a21oi_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _07223_ _07224_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__xnor2_1
X_11663_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04808_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__and3_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13402_ _06069_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10614_ _03908_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14382_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _07144_ VGND
+ VGND VPWR VPWR _07166_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11594_ _03619_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13333_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _06247_ VGND VGND
+ VPWR VPWR _06262_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10545_ _03535_ _03846_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13264_ _06202_ net148 _06203_ _06206_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10476_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03773_ _03651_
+ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__o21ai_1
X_15003_ clknet_leaf_107_i_clk _00548_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12215_ _05292_ _05293_ _05296_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13195_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06142_ _06138_
+ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12146_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or4_4
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05172_
+ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__or2_1
X_11028_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _04251_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12979_ _05954_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14718_ clknet_leaf_53_i_clk _00263_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14649_ clknet_leaf_49_i_clk _00194_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08170_ _01703_ _01758_ _01759_ _01730_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_7_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR out_sintheta[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07954_ _01557_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__xor2_2
X_07885_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\] _01499_ _01480_ VGND
+ VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09624_ _02595_ _03038_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09555_ _02975_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08506_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR VPWR
+ _02047_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09486_ _02905_ _02908_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08437_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\] _01983_ VGND VGND VPWR
+ VPWR _01984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08368_ _01891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _01923_ _01925_ _01908_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07319_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _01045_ _01062_
+ _01064_ _01059_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08299_ _01868_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10330_ _03654_ _03652_ _03653_ _03631_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10261_ _03603_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__clkbuf_1
X_12000_ _05115_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__and2_1
X_10192_ _03539_ _03542_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13951_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06795_ VGND
+ VGND VPWR VPWR _06796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12902_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _05885_
+ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__or2_1
X_13882_ _06734_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__nand2_1
X_12833_ _05835_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _05774_ _05775_ _05489_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__o21ai_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _04754_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__clkbuf_4
X_14503_ clknet_leaf_4_i_clk _00049_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05711_ VGND
+ VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xnor2_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11646_ _04802_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14434_ _07209_ _07204_ _07206_ _01861_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__o31a_1
Xinput14 in_alpha[3] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_0_80_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14365_ _07059_ _07150_ _07151_ _01475_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 in_x[13] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
X_11577_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _04723_ VGND
+ VGND VPWR VPWR _04750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput36 in_x[7] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xinput47 in_y[17] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
X_13316_ _05927_ _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10528_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__and2b_1
X_14296_ _07081_ _07090_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13247_ _06192_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10459_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03770_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13178_ _06115_ _06124_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__or2b_1
X_12129_ _05217_ _05219_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07670_ net15 net16 net17 VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__or3_2
X_09340_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _02783_
+ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09271_ _02715_ _02723_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08222_ _01803_ _01804_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08153_ _01472_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08084_ net41 net23 VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08986_ _02471_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _02472_ sky130_fd_sc_hd__or2b_1
X_07937_ _01543_ _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__or2b_1
X_07868_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[5\] _01484_
+ _01486_ _01475_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09607_ _02754_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _03017_
+ _03023_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__o211a_1
X_07799_ net4 _01431_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__nand2_1
X_09538_ _02957_ _02958_ _02960_ _02928_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__a221o_2
XFILLER_0_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09469_ _02893_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11500_ _04444_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _04682_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12480_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__clkbuf_4
X_11431_ _04468_ _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14150_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR _06966_ sky130_fd_sc_hd__inv_2
X_11362_ _04549_ _04553_ _04547_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13101_ _05854_ net314 _05847_ _06062_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03640_
+ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__and2_1
X_14081_ _06905_ net263 _06678_ _06908_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11293_ _04444_ net479 VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__or2_1
X_13032_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _06003_ VGND
+ VGND VPWR VPWR _06004_ sky130_fd_sc_hd__xnor2_1
X_10244_ _03190_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND
+ VGND VPWR VPWR _03590_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10175_ _03190_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _03528_ sky130_fd_sc_hd__or2_1
X_14983_ clknet_leaf_95_i_clk _00528_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13934_ _06779_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__nor2_1
X_13865_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ _06707_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12816_ _05819_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13796_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _06660_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12747_ _05755_ _05758_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__and2_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12678_ _05652_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11629_ _04773_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _04785_ _04787_ _04788_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14417_ _07172_ _07194_ _07195_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15397_ clknet_leaf_30_i_clk _00942_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14348_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _07133_ _07135_
+ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14279_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _07023_ VGND
+ VGND VPWR VPWR _07076_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _02340_ _02345_ net469 VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _02286_ _02287_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__nor2_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_3_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_07722_ _01379_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_100_i_clk clknet_4_4_0_i_clk VGND VGND VPWR VPWR clknet_leaf_100_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07653_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] VGND VGND VPWR VPWR
+ _01328_ sky130_fd_sc_hd__inv_2
X_07584_ _01271_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_115_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_115_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09323_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _02773_
+ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09254_ _02711_ _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08205_ _01577_ _01584_ _01789_ _01576_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09185_ _02608_ _02627_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__or3_1
X_08136_ _01691_ _01706_ _01707_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08067_ net22 net40 VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08969_ _02321_ net619 _02381_ _02456_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__o211a_1
X_11980_ _05098_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__xor2_1
X_10931_ _04048_ _04182_ _04183_ _04063_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10862_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04119_ VGND
+ VGND VPWR VPWR _04120_ sky130_fd_sc_hd__xor2_1
X_13650_ _06516_ _06523_ _06529_ _06536_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _05619_ _05623_ _05629_ _05487_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__a31o_1
X_13581_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _06463_ VGND
+ VGND VPWR VPWR _06479_ sky130_fd_sc_hd__or2_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _04023_ net422 _04057_ _04058_ _04059_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__o221a_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR
+ VPWR _05569_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15320_ clknet_leaf_18_i_clk _00865_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12463_ _05500_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _05510_ _05511_ _05391_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__o221a_1
X_15251_ clknet_leaf_5_i_clk _00796_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_11414_ _04390_ net331 _04387_ _04603_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14202_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _07007_ VGND
+ VGND VPWR VPWR _07009_ sky130_fd_sc_hd__and2_1
X_15182_ clknet_leaf_115_i_clk _00727_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12394_ _05450_ _05453_ _05452_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14133_ _06646_ _06951_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__nand2_1
X_11345_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ _04518_ _04542_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__o31a_1
XFILLER_0_151_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14064_ _06865_ _06894_ _06890_ _06891_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11276_ _04478_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13015_ _05986_ _05987_ _05841_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__a21o_1
X_10227_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__inv_2
X_10158_ _03498_ _03503_ _03497_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14966_ clknet_leaf_95_i_clk _00511_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_10089_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__and2b_1
X_13917_ _06761_ _06766_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__xor2_1
X_14897_ clknet_leaf_87_i_clk _00442_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_32_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13848_ _06561_ net599 _06678_ _06706_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13779_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _06646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold403 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND VGND VPWR
+ VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold414 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net531 sky130_fd_sc_hd__buf_1
Xhold425 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR VPWR
+ net542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold436 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold447 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND VGND VPWR
+ VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold458 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] VGND VGND VPWR
+ VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _03205_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03255_
+ _03183_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _02324_
+ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__nand2_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _02257_ _02271_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__nand2_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _01338_ _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__nand2_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _01880_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[13\] _01314_ _01282_
+ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07567_ net206 _01260_ _01255_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09306_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07498_ _01016_ net231 _01216_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09237_ _02698_ _02694_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09168_ _02497_ _02636_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08119_ _01709_ _01711_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09099_ _02564_ _02568_ _02573_ _02369_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11130_ _04336_ _04350_ _04351_ _04357_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__and4_1
X_11061_ _04298_ _04299_ _03994_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a21o_1
X_10012_ _03201_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03379_
+ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__a22o_1
X_14820_ clknet_leaf_110_i_clk net146 VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14751_ clknet_leaf_65_i_clk _00296_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_11963_ _05084_ _05085_ _04786_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__o21ai_1
X_13702_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _06571_
+ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__nand2_1
X_10914_ _04166_ _04167_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__a21o_1
X_11894_ _05021_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__and2b_1
X_14682_ clknet_leaf_62_i_clk _00227_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10845_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _04095_ _04097_
+ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13633_ _06515_ _06522_ _06523_ _06200_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10776_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04044_
+ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__xnor2_1
X_13564_ _06461_ _06463_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15303_ clknet_leaf_13_i_clk _00848_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12515_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05550_
+ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13495_ _06403_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12446_ _05490_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__or2_1
X_15234_ clknet_leaf_14_i_clk _00779_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12377_ _05222_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05441_
+ _05442_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15165_ clknet_leaf_110_i_clk net154 VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11328_ _04523_ _04526_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__or3_1
X_14116_ _06935_ _06936_ _06937_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__a21oi_1
X_15096_ clknet_leaf_117_i_clk _00641_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11259_ _04457_ _04458_ _04463_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__o31a_1
X_14047_ _06878_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__xnor2_1
X_14949_ clknet_leaf_106_i_clk _00494_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_08470_ _02013_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07421_ _01154_ _01155_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07352_ _01044_ net185 _01094_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07283_ _01016_ net243 _01028_ _01031_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09022_ _02343_ _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold200 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 net91 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold244 diff3\[16\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 net59 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold266 diff3\[12\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 diff2\[12\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 net84 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _03293_ _03294_ _03299_ _03185_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _03237_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _03241_ _03242_ _03013_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__o221a_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _02314_ net191 _01945_ _02317_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09786_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _03185_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _02217_ _02253_ _02254_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__a211o_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[6\] _02193_ VGND VGND VPWR
+ VPWR _02194_ sky130_fd_sc_hd__xnor2_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ diff2\[10\] _01270_ _01272_ diff3\[10\] _01300_ VGND VGND VPWR VPWR _01301_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _02118_ _02131_ _02132_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10630_ _03708_ _03922_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10561_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _03861_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12300_ _05372_ _03118_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13280_ _06210_ net598 _06215_ _06217_ _06197_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10492_ _03626_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03798_
+ _03800_ _03633_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__o221a_1
XFILLER_0_106_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12231_ _05234_ _05311_ _05312_ _05080_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12162_ _05248_ _05249_ _01250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11113_ _04339_ _04341_ _04345_ _04047_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12093_ _05153_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _05189_ _05190_ _05170_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__o221a_1
X_11044_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04283_ VGND
+ VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14803_ clknet_leaf_74_i_clk _00348_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12995_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05969_ VGND
+ VGND VPWR VPWR _05970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14734_ clknet_leaf_71_i_clk _00279_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11946_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05069_
+ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__nor2_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14665_ clknet_leaf_54_i_clk _00210_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11877_ _05005_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13616_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _06488_ VGND
+ VGND VPWR VPWR _06510_ sky130_fd_sc_hd__xor2_1
X_10828_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04089_ _03996_
+ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__mux2_1
X_14596_ clknet_leaf_46_i_clk _00141_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13547_ _06069_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__and2_1
X_10759_ _04028_ _04029_ _03669_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13478_ _06383_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15217_ clknet_leaf_2_i_clk _00762_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12429_ _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15148_ clknet_leaf_121_i_clk _00693_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07970_ _01565_ _01571_ _01573_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__o21ai_1
X_15079_ clknet_leaf_119_i_clk _00624_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_09640_ _03039_ _03043_ _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09571_ _02992_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
X_08522_ _01998_ _02005_ _02014_ _02030_ _02041_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08453_ _01984_ _01991_ _01997_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07404_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _01051_ _01052_
+ _01140_ _01057_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08384_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] _01932_ _01549_
+ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07335_ _01077_ _01078_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07266_ _01012_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09005_ _02481_ _02488_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09907_ _03237_ net431 _03284_ _03285_ _03258_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__o221a_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _03221_
+ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__and2_1
X_09769_ _03162_ _03163_ _03164_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__o21ba_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _04925_ _04936_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__nor2_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _05789_ _05783_
+ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__a21oi_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11731_ _04875_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__and2b_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _07157_ VGND
+ VGND VPWR VPWR _07224_ sky130_fd_sc_hd__xnor2_1
X_11662_ _04773_ net566 _04815_ _04816_ _04788_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13401_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _06320_ _06204_
+ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__mux2_1
X_10613_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03907_ VGND
+ VGND VPWR VPWR _03909_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11593_ _04756_ net122 _04387_ _04761_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__o211a_1
X_14381_ _07165_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10544_ _03605_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _03844_
+ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__a22o_1
X_13332_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _06260_ _06261_ _06197_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10475_ _03768_ _03781_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__or2_1
X_13263_ net647 _06205_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15002_ clknet_leaf_107_i_clk _00547_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12214_ _01249_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13194_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _06142_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12145_ _05228_ _05230_ _05227_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12076_ _05140_ net643 _05141_ _05176_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__o211a_1
X_11027_ _04023_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _04267_
+ _04268_ _04059_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__o221a_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12978_ _05944_ _05946_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14717_ clknet_leaf_53_i_clk _00262_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11929_ _04771_ net533 _05053_ _05054_ _04965_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14648_ clknet_leaf_32_i_clk _00193_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14579_ clknet_leaf_40_i_clk _00124_ VGND VGND VPWR VPWR diff3\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput102 net102 VGND VGND VPWR VPWR out_sintheta[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07953_ net21 net39 VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07884_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\] _01499_ VGND VGND
+ VPWR VPWR _01500_ sky130_fd_sc_hd__nor2_1
X_09623_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03037_ VGND
+ VGND VPWR VPWR _03038_ sky130_fd_sc_hd__xnor2_1
X_09554_ _02962_ _02976_ _02967_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__a21bo_1
X_08505_ _01867_ _02045_ _02046_ _01552_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09485_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _02913_ VGND
+ VGND VPWR VPWR _02914_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08436_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[4\] _01982_ VGND VGND VPWR
+ VPWR _01983_ sky130_fd_sc_hd__xnor2_1
X_08367_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[10\] _01921_ _01922_
+ _01924_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07318_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _01051_ _01052_
+ _01063_ _01057_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a221o_1
X_08298_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_out VGND VGND VPWR VPWR _01868_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07249_ _01004_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10260_ _03186_ _02310_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10191_ _03519_ _03526_ _03531_ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13950_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06587_ VGND VGND
+ VPWR VPWR _06795_ sky130_fd_sc_hd__o31a_1
X_12901_ _05854_ net575 _05847_ _05889_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__o211a_1
X_13881_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06684_ VGND
+ VGND VPWR VPWR _06735_ sky130_fd_sc_hd__or2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _05652_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__and2_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12763_ _05759_ _05762_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__or2b_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14502_ clknet_leaf_4_i_clk _00048_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _04861_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12694_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _05525_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__o21a_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _07204_ _07206_ _07209_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__o21ai_1
X_11645_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _04789_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14364_ _06909_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _07151_ sky130_fd_sc_hd__or2_1
Xinput15 in_alpha[4] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
X_11576_ _04742_ _04745_ _04741_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 in_x[14] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 in_x[8] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput48 in_y[1] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
X_13315_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06242_
+ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__or2_1
X_10527_ _03625_ net455 _03620_ _03830_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__o211a_1
X_14295_ _07078_ _07084_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__nor2_1
X_13246_ _06069_ _06191_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__and2_1
X_10458_ _03765_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13177_ _06126_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__inv_2
X_10389_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND
+ VGND VPWR VPWR _03707_ sky130_fd_sc_hd__or2_1
X_12128_ _05217_ _05219_ _05128_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__a21o_1
X_12059_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _05160_
+ _01250_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09270_ _02728_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08221_ _01529_ net508 _01794_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08152_ _01738_ _01742_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08083_ _01463_ net514 _01635_ _01678_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08985_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _02470_ VGND
+ VGND VPWR VPWR _02471_ sky130_fd_sc_hd__xor2_1
X_07936_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[15\]
+ _01534_ _01328_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__a31o_1
X_07867_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[5\] _01483_ _01485_ VGND
+ VGND VPWR VPWR _01486_ sky130_fd_sc_hd__o21ai_1
X_09606_ _03021_ _03022_ _02755_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07798_ _01431_ _01432_ net248 _01333_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__o2bb2a_1
X_09537_ _02944_ _02959_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09468_ _02888_ _02897_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08419_ _01873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _01968_ sky130_fd_sc_hd__or2_1
X_09399_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _02837_
+ _02751_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11430_ _04375_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _04616_
+ _04617_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11361_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04545_ VGND
+ VGND VPWR VPWR _04558_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13100_ _06060_ _06061_ _05855_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__o21ai_1
X_10312_ _03280_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _03629_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__o31a_1
X_11292_ _04493_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__xnor2_1
X_14080_ _06907_ _01022_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13031_ _05982_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__buf_4
X_10243_ _03587_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__xnor2_1
X_10174_ _03519_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__xor2_1
X_14982_ clknet_leaf_95_i_clk _00527_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_13933_ _06778_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _06780_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13864_ _06556_ _06719_ _06720_ _06459_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__o211a_1
X_12815_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05789_ VGND
+ VGND VPWR VPWR _05820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13795_ _06651_ _06655_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12746_ _05755_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _05486_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05696_
+ _05697_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14416_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _07157_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__o41a_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11628_ _04538_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__clkbuf_4
X_15396_ clknet_leaf_30_i_clk _00941_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ _07134_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR VPWR
+ _07135_ sky130_fd_sc_hd__mux2_1
X_11559_ _04727_ _04734_ _02132_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14278_ _06905_ _07074_ _07075_ _06996_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13229_ _06175_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__and2b_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _02275_ _02278_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__nand2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07721_ _01378_ net445 _01344_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07652_ _01327_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
X_07583_ diff2\[17\] _01259_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09322_ _02763_ _02768_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09253_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _02713_ VGND
+ VGND VPWR VPWR _02714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08204_ _01565_ _01780_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09184_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08135_ _01722_ _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08066_ net40 net22 VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08968_ _02453_ _02454_ _02455_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__o21ai_1
X_07919_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[13\] _01526_ _01527_
+ _01529_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__o31ai_1
X_08899_ _02393_ _02395_ _02344_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__mux2_1
X_10930_ _04010_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _04183_ sky130_fd_sc_hd__or2_1
X_10861_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04108_ _04034_
+ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12600_ _05619_ _05623_ _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__a21oi_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13580_ _06478_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10792_ _02308_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _05488_ _05565_ _05568_ _05343_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__o211a_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15250_ clknet_4_2_0_i_clk _00795_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12462_ _05505_ _05509_ _05487_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14201_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _07007_ VGND
+ VGND VPWR VPWR _07008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11413_ _04601_ _04602_ _04391_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15181_ clknet_leaf_115_i_clk _00726_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12393_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05423_ VGND
+ VGND VPWR VPWR _05456_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14132_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _06940_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__and3_1
X_11344_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR _04542_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14063_ _06865_ _06890_ _06891_ _06894_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__o31ai_2
X_11275_ _04462_ _04464_ _04473_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a21boi_2
X_13014_ _05986_ _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__nor2_1
X_10226_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03572_ _03573_
+ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__or3_2
X_10157_ _03509_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__or2_1
X_14965_ clknet_leaf_89_i_clk _00510_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_4
X_10088_ _03189_ net297 _03017_ _03448_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__o211a_1
X_13916_ _06739_ _06763_ _06765_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__and3_1
X_14896_ clknet_leaf_106_i_clk _00441_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_13847_ _06563_ _06705_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13778_ _06563_ net442 _06644_ _06645_ _06631_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12729_ _05632_ _05742_ _05743_ _05675_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15379_ clknet_leaf_38_i_clk _00924_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
Xmax_cap112 net113 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xhold404 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR
+ VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold415 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND VGND VPWR
+ VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND VGND VPWR
+ VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09940_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__or4_4
Xhold459 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _03255_
+ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__nor2_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _02324_
+ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__or2_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _02252_ _02263_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07704_ net7 _01361_ net8 VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__a21o_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\]
+ _02170_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__or4_4
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ r_i_alpha1\[13\] _01313_ _01258_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__mux2_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09305_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07497_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _01159_ _01214_
+ _01215_ _01030_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09236_ _02694_ _02698_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09167_ _02319_ _02631_ _02633_ _02635_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08118_ _01691_ _01697_ _01710_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09098_ _02564_ _02568_ _02573_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08049_ _01625_ _01646_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11060_ _04291_ _04297_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10011_ _03373_ _03378_ _03185_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14750_ clknet_leaf_65_i_clk _00295_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11962_ _05082_ _05083_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__and2_1
X_13701_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _06567_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__or3_1
X_10913_ _04164_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04150_
+ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__or3_1
X_14681_ clknet_leaf_63_i_clk _00226_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11893_ _05013_ _05020_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__nand2_1
X_13632_ _06515_ _06522_ _06523_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__a21oi_1
X_10844_ _04102_ _04103_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13563_ _06462_ _05927_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__mux2_2
XFILLER_0_82_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10775_ _04041_ _04043_ _04035_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15302_ clknet_leaf_13_i_clk _00847_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12514_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _05553_ _05554_ _05544_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13494_ _06069_ _06402_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15233_ clknet_leaf_14_i_clk net558 VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12445_ _05488_ net269 _05495_ _05497_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15164_ clknet_leaf_110_i_clk net150 VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12376_ _05439_ _05440_ _01249_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR _06937_ sky130_fd_sc_hd__inv_2
X_11327_ _04478_ _04479_ _04505_ _04497_ _04514_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__o2111a_1
X_15095_ clknet_leaf_118_i_clk _00640_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046_ _06866_ _06879_ _06871_ _06862_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__o211a_1
X_11258_ _04457_ _04458_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_114_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_114_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_157_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10209_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND VGND VPWR
+ VPWR _03558_ sky130_fd_sc_hd__inv_2
X_11189_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _04404_
+ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__and2_1
X_14948_ clknet_leaf_106_i_clk _00493_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14879_ clknet_leaf_110_i_clk net142 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07420_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _01146_ VGND
+ VGND VPWR VPWR _01155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07351_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _01045_ _01091_
+ _01093_ _01059_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07282_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _01029_ _01030_
+ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09021_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ _02483_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold201 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net318 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold212 r_i_alpha1\[9\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold223 diff1\[12\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _00713_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 diff1\[15\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold256 net70 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 net74 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _03293_ _03294_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold289 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ net603 _03240_ _03183_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__a21o_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _02315_
+ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__or2_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _03183_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08736_ _02241_ _02255_ _02245_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__a21oi_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08667_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[7\] _02192_ VGND VGND VPWR
+ VPWR _02193_ sky130_fd_sc_hd__xnor2_2
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_i_clk clknet_4_5_0_i_clk VGND VGND VPWR VPWR clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _01273_ diff1\[10\] VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__and2_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _01794_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07549_ net65 net432 _01012_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10560_ _03852_ _03854_ _03859_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09219_ _02669_ _02683_ _02132_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10491_ _03642_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12230_ _05139_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _05312_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12161_ _05248_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_31_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11112_ _04339_ _04341_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12092_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05188_
+ _05129_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__a21o_1
X_11043_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04282_ VGND
+ VGND VPWR VPWR _04283_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_46_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14802_ clknet_leaf_74_i_clk _00347_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_12994_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05961_ _05877_
+ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14733_ clknet_leaf_72_i_clk _00278_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_11945_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05059_ VGND
+ VGND VPWR VPWR _05069_ sky130_fd_sc_hd__nor2_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ clknet_leaf_58_i_clk _00209_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11876_ _05002_ _05004_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13615_ _06505_ _06504_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10827_ _04087_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14595_ clknet_leaf_46_i_clk _00140_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13546_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _06447_ _06204_
+ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux2_1
X_10758_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04018_
+ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13477_ _06385_ _06387_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__and2_1
X_10689_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03944_ VGND
+ VGND VPWR VPWR _03977_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15216_ clknet_leaf_2_i_clk _00761_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12428_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05485_ sky130_fd_sc_hd__inv_2
X_15147_ clknet_leaf_125_i_clk _00692_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12359_ _05425_ _05416_ _05419_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15078_ clknet_leaf_120_i_clk _00623_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14029_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _06845_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__o41a_1
X_09570_ _02497_ _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08521_ _02059_ _02060_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08452_ _01984_ _01991_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_148_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07403_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _01132_ VGND
+ VGND VPWR VPWR _01140_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08383_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[11\]
+ _01928_ _01549_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07334_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _01066_ VGND
+ VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07265_ _01014_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09004_ _02481_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09906_ _03283_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _03183_
+ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _03207_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__or2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _03138_ _03156_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__and3_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _02240_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09699_ _03048_ _03068_ _03086_ _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__or4_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _04874_ VGND
+ VGND VPWR VPWR _04876_ sky130_fd_sc_hd__or2b_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11661_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04814_
+ _04786_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__o21ai_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13400_ _06318_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__xor2_1
X_10612_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03907_ VGND
+ VGND VPWR VPWR _03908_ sky130_fd_sc_hd__nand2_1
X_14380_ _01253_ _07164_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__and2_1
X_11592_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] _04758_
+ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13331_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _06259_
+ _06201_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10543_ _03841_ _03843_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13262_ _06204_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__buf_2
X_10474_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03775_ _03783_
+ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_122_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15001_ clknet_leaf_107_i_clk _00546_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12213_ _05292_ _05293_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__or3b_1
XFILLER_0_121_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13193_ _05998_ _06144_ _06145_ _06110_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12144_ _05222_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12075_ _05142_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__nand2_1
X_11026_ _04254_ _04259_ _04266_ _03994_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12977_ _05952_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11928_ _05036_ _05045_ _05052_ _04755_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__a31o_1
X_14716_ clknet_leaf_53_i_clk _00261_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14647_ clknet_leaf_44_i_clk _00192_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_11859_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _04990_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14578_ clknet_leaf_39_i_clk _00123_ VGND VGND VPWR VPWR diff1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13529_ _06232_ _06431_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput103 net103 VGND VGND VPWR VPWR out_sintheta[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07952_ net30 net48 VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__xor2_4
X_07883_ _01497_ _01498_ _01329_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__mux2_1
X_09622_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02769_ VGND VGND VPWR
+ VPWR _03037_ sky130_fd_sc_hd__o31a_1
X_09553_ _02969_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__inv_2
X_08504_ _01873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _02046_ sky130_fd_sc_hd__or2_1
X_09484_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _02912_ VGND
+ VGND VPWR VPWR _02913_ sky130_fd_sc_hd__xor2_2
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08435_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[3\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\] _01879_ VGND VGND VPWR VPWR
+ _01982_ sky130_fd_sc_hd__o31a_1
X_08366_ _01865_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07317_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _01053_ VGND
+ VGND VPWR VPWR _01063_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08297_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__buf_4
XFILLER_0_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07248_ net367 _01003_ _01000_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10190_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03530_ _03540_
+ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__o21ai_1
X_12900_ _05855_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__nand2_1
X_13880_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06684_ VGND
+ VGND VPWR VPWR _06734_ sky130_fd_sc_hd__nand2_1
X_12831_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05833_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _05772_ _05773_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__or2_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14501_ clknet_leaf_4_i_clk _00047_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _04850_ _04860_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__and2_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _05632_ _05709_ _05710_ _05675_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__o211a_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _07207_ _07208_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__and2_1
X_11644_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _04778_ VGND VGND
+ VPWR VPWR _04801_ sky130_fd_sc_hd__and4_1
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14363_ _07148_ _07149_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11575_ _04748_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
Xinput16 in_alpha[5] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput27 in_x[15] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
X_13314_ _06210_ net637 _06203_ _06246_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__o211a_1
Xinput38 in_x[9] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
X_10526_ _03828_ _03829_ _03642_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_135_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 in_y[2] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
X_14294_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _07041_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13245_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06190_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__mux2_1
X_10457_ _03743_ _03766_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13176_ _06106_ _06103_ _06104_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__o21ba_1
X_10388_ _03699_ _03705_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__xnor2_1
X_12127_ _05206_ _05210_ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__o21a_1
X_12058_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _05160_
+ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__and2_1
X_11009_ _04034_ _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08220_ _01572_ _01621_ _01801_ _01802_ _01457_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08151_ _01722_ _01726_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08082_ _01562_ _01667_ _01677_ _01485_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08984_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _02442_ _02341_ VGND
+ VGND VPWR VPWR _02470_ sky130_fd_sc_hd__o41a_1
X_07935_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[15\]
+ _01531_ _01328_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__o31a_1
X_07866_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in VGND VGND VPWR VPWR _01485_
+ sky130_fd_sc_hd__buf_4
X_09605_ _03014_ _03020_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07797_ net20 _01428_ _01344_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09536_ _02940_ _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09467_ _02894_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08418_ _01962_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09398_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _02837_
+ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08349_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND VPWR VPWR
+ _01909_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11360_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR
+ VPWR _04557_ sky130_fd_sc_hd__clkbuf_4
X_10311_ _03280_ _03634_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11291_ _04480_ _04486_ _04484_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13030_ _05952_ _05959_ _05986_ _06001_ _05994_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__a2111o_1
X_10242_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03572_ VGND
+ VGND VPWR VPWR _03588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_784 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10173_ _03524_ _03525_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14981_ clknet_leaf_89_i_clk _00526_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_13932_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _06778_ VGND
+ VGND VPWR VPWR _06779_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13863_ _06557_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND
+ VGND VPWR VPWR _06720_ sky130_fd_sc_hd__or2_1
X_12814_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05789_ VGND
+ VGND VPWR VPWR _05819_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13794_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _06654_ VGND
+ VGND VPWR VPWR _06658_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12745_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05757_ VGND
+ VGND VPWR VPWR _05758_ sky130_fd_sc_hd__xnor2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _05670_ _05695_ _05691_ _05692_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__o41a_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14415_ _07175_ _07183_ _07188_ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__and3_1
X_11627_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _04784_
+ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15395_ clknet_leaf_30_i_clk _00940_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14346_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _07133_
+ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__nor2_1
X_11558_ _04732_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10509_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03796_ VGND
+ VGND VPWR VPWR _03815_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14277_ _06907_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND
+ VGND VPWR VPWR _07075_ sky130_fd_sc_hd__or2_1
X_11489_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ _04632_ _04670_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__or4_4
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13228_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06136_ VGND
+ VGND VPWR VPWR _06176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06114_ VGND
+ VGND VPWR VPWR _06115_ sky130_fd_sc_hd__and2_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _00991_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07651_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[16\] _01326_ diff_valid
+ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07582_ _01269_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09321_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__buf_4
X_09252_ _01958_ _02712_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08203_ _01717_ net631 _01635_ _01788_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09183_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR _02650_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08134_ _01724_ _01725_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08065_ _01539_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\] _01657_ _01660_
+ _01661_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08967_ _02453_ _02454_ _02333_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__a21oi_1
X_07918_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in VGND VGND VPWR VPWR _01529_
+ sky130_fd_sc_hd__buf_4
X_08898_ _02394_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__inv_2
X_07849_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] VGND VGND VPWR VPWR
+ _01470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10860_ _04118_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09519_ _02928_ _02941_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__a21bo_1
X_10791_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _04056_
+ _03994_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _05492_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ _05505_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14200_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _07006_ VGND
+ VGND VPWR VPWR _07007_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11412_ net282 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _04602_ sky130_fd_sc_hd__nor2_1
X_15180_ clknet_leaf_115_i_clk _00725_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12392_ _05234_ _05454_ _05455_ _05343_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__o211a_1
X_14131_ _06905_ _06949_ _06950_ _06747_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11343_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ _04518_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__nor3_1
XFILLER_0_1_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14062_ _06892_ _06893_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11274_ _04471_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13013_ _05972_ _05975_ _05971_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__a21oi_1
X_10225_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03569_ VGND
+ VGND VPWR VPWR _03573_ sky130_fd_sc_hd__and2_1
X_10156_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03508_ VGND
+ VGND VPWR VPWR _03510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
X_14964_ clknet_leaf_93_i_clk _00509_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_10087_ _03446_ _03447_ _03191_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__o21ai_1
X_13915_ _06749_ _06764_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__nor2_1
X_14895_ clknet_leaf_81_i_clk _00440_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13846_ _06703_ _06704_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13777_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _06642_
+ _06643_ _06584_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__o31ai_1
X_10989_ _03996_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12728_ _05499_ net641 VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12659_ _05669_ _05670_ _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15378_ clknet_leaf_29_i_clk _00923_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold405 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ _07113_ _07118_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__or2_1
Xhold416 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold427 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND VGND VPWR
+ VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold438 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR VPWR
+ net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09870_ _03249_ _03253_ _02850_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__mux2_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _02315_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__clkbuf_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\] _02262_ _02269_ VGND
+ VGND VPWR VPWR _02270_ sky130_fd_sc_hd__o21ai_2
X_07703_ net7 net8 _01361_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__and3_1
X_08683_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[7\]
+ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07634_ diff2\[13\] _01270_ _01272_ diff3\[13\] _01312_ VGND VGND VPWR VPWR _01313_
+ sky130_fd_sc_hd__a221o_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07565_ _01257_ diff2\[17\] _01258_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_137_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09304_ _02750_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07496_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _01122_ _01140_
+ _01046_ _01072_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09235_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _02697_ VGND
+ VGND VPWR VPWR _02698_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09166_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out _02634_ VGND
+ VGND VPWR VPWR _02635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08117_ net24 net42 VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09097_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _02555_ VGND
+ VGND VPWR VPWR _02573_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08048_ _01614_ _01615_ _01644_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10010_ _03373_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nand2_1
X_09999_ _03359_ _03364_ _03367_ _03201_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a31o_1
X_11961_ _05082_ _05083_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10912_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ _04165_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__a21oi_2
X_13700_ _06565_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _06578_ _06579_ _06526_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__o221a_1
X_14680_ clknet_leaf_63_i_clk _00225_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_11892_ _05013_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13631_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06514_ VGND
+ VGND VPWR VPWR _06523_ sky130_fd_sc_hd__xor2_2
X_10843_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _04101_ VGND
+ VGND VPWR VPWR _04103_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13562_ _05927_ _06460_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10774_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12513_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05552_
+ _05490_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__o21ai_1
X_15301_ clknet_leaf_18_i_clk _00846_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13493_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06401_ _06204_
+ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15232_ clknet_leaf_12_i_clk _00777_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12444_ net176 _05492_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15163_ clknet_leaf_15_i_clk _00708_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12375_ _05439_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ _06917_ _06934_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__a31o_1
X_11326_ _04505_ _04499_ _04514_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__a31o_1
X_15094_ clknet_leaf_120_i_clk _00639_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14045_ _06863_ _06872_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__nand2_1
X_11257_ _04461_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10208_ _03539_ _03541_ _03548_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__or3_1
X_11188_ _04061_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _04394_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__o31a_1
X_10139_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _03494_ sky130_fd_sc_hd__inv_2
X_14947_ clknet_leaf_106_i_clk _00492_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14878_ clknet_leaf_110_i_clk net133 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13829_ _06561_ net639 _06678_ _06690_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07350_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _01051_ _01052_
+ _01092_ _01057_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07281_ _01012_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09020_ _02481_ _02502_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold202 _01231_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold213 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 r_i_alpha1\[7\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND VGND VPWR
+ VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 r_i_alpha1\[14\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 net88 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 net94 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09922_ _03297_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__and2_1
Xhold279 diff3\[15\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09853_ net580 _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__nor2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _02314_ net155 _01945_ _02316_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__o211a_1
X_09784_ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__clkbuf_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\] _02243_ VGND VGND VPWR
+ VPWR _02255_ sky130_fd_sc_hd__nand2_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _01880_ _02191_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__and2_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07617_ _01299_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _02129_ _02130_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__nor2_1
X_07548_ _01246_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07479_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _01081_ _01085_
+ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09218_ _02681_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10490_ _03789_ _03792_ _03797_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__or3b_1
X_09149_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _02618_ VGND
+ VGND VPWR VPWR _02619_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ _05235_ _05241_ _05239_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11111_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04338_ VGND
+ VGND VPWR VPWR _04345_ sky130_fd_sc_hd__xor2_1
X_12091_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05188_
+ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11042_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _04281_ _04035_
+ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14801_ clknet_leaf_74_i_clk _00346_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12993_ _05843_ _05967_ _05968_ _05938_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__o211a_1
X_14732_ clknet_leaf_72_i_clk _00277_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_11944_ _04862_ _05067_ _05068_ _04739_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11875_ _05002_ _05004_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__nor2_1
X_14663_ clknet_leaf_54_i_clk _00208_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10826_ _04077_ _04079_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__nand2_1
X_13614_ _06508_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14594_ clknet_leaf_49_i_clk _00139_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10757_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _04015_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__or3_1
X_13545_ _06445_ _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13476_ _06374_ _06386_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10688_ _01765_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15215_ clknet_leaf_124_i_clk _00760_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_113_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12427_ _05484_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12358_ _05416_ _05419_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__a21oi_1
X_15146_ clknet_leaf_121_i_clk _00691_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11309_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04500_ _04413_
+ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15077_ clknet_leaf_119_i_clk _00622_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_12289_ _05362_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14028_ _06844_ _06851_ _06858_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__and3_1
X_08520_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[10\] _02058_ VGND VGND VPWR
+ VPWR _02060_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08451_ _01995_ _01996_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07402_ _01019_ _01138_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08382_ _01891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _01936_ _01937_ _01908_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07333_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _01066_ VGND
+ VGND VPWR VPWR _01077_ sky130_fd_sc_hd__or2_4
XFILLER_0_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07264_ net385 _01011_ _01013_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09003_ _02486_ _02487_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09905_ _03283_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _03284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _03216_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__or3_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _03153_ _03165_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__nor2_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _01981_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__and2_1
X_09698_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__or2_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _02161_ _02165_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__o21a_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04814_
+ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__and2_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_113_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_113_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10611_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03906_ VGND
+ VGND VPWR VPWR _03907_ sky130_fd_sc_hd__xnor2_1
X_11591_ _04756_ net128 _04387_ _04760_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13330_ net483 _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10542_ _03841_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13261_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _06204_ sky130_fd_sc_hd__clkbuf_4
X_10473_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03775_ _03763_
+ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12212_ _05294_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__or2_1
X_15000_ clknet_leaf_107_i_clk net286 VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13192_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _06145_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12143_ _05233_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12074_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05174_
+ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__xnor2_1
X_11025_ _04254_ _04259_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12976_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05951_ VGND
+ VGND VPWR VPWR _05953_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14715_ clknet_leaf_53_i_clk _00260_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11927_ _05036_ _05045_ _05052_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14646_ clknet_leaf_43_i_clk _00191_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _04984_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _04989_ sky130_fd_sc_hd__and2b_1
XFILLER_0_68_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10809_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _04068_ VGND
+ VGND VPWR VPWR _04072_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11789_ _04862_ _04928_ _04929_ _04739_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__o211a_1
X_14577_ clknet_leaf_42_i_clk _00122_ VGND VGND VPWR VPWR diff1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13528_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _06431_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13459_ _06201_ net409 VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput104 net104 VGND VGND VPWR VPWR out_sintheta[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15129_ clknet_leaf_122_i_clk _00674_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_i_clk clknet_4_5_0_i_clk VGND VGND VPWR VPWR clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07951_ _01470_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07882_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] _01489_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[7\]
+ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09621_ _02591_ _03027_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__or2_1
X_09552_ _02972_ _02974_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__xnor2_1
X_08503_ _02043_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__and2_1
X_09483_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _02902_ _02770_
+ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_i_clk clknet_4_10_0_i_clk VGND VGND VPWR VPWR clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08434_ _01765_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08365_ _01921_ _01922_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[10\]
+ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07316_ _01019_ _01061_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08296_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_45_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07247_ net6 VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09819_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _03198_
+ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12830_ _05829_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__xor2_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _05768_ _05771_
+ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__nor3_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ clknet_leaf_25_i_clk _00046_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _04857_ _04859_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ _04754_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _05499_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _05710_ sky130_fd_sc_hd__or2_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _04773_ net625 _04799_ _04800_ _04788_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__o221a_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14431_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _07156_ VGND
+ VGND VPWR VPWR _07208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11574_ _04468_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__and2_4
X_14362_ _07143_ _07139_ _07147_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 in_alpha[6] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 in_x[16] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
X_10525_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__nor2_1
X_13313_ _06232_ _06245_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__nand2_1
Xinput39 in_y[0] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_0_80_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14293_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _07041_ VGND
+ VGND VPWR VPWR _07088_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13244_ _06186_ _06189_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10456_ _03752_ _03754_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13175_ _05855_ net388 _06127_ _06129_ _05910_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__o221a_1
X_10387_ _03703_ _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12126_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _05209_ VGND
+ VGND VPWR VPWR _05218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12057_ _05158_ _05159_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11008_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__or4_2
XFILLER_0_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12959_ _04455_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14629_ clknet_leaf_44_i_clk _00174_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_08150_ net26 net44 VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08081_ _01669_ _01675_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08983_ _02469_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07934_ _01539_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[15\] _01541_
+ _01542_ _01513_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__o221a_1
X_07865_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[5\] _01483_ VGND VGND
+ VPWR VPWR _01484_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _03014_ _03020_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07796_ net20 _01428_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09535_ _02939_ _02953_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09466_ _02844_ net585 _02895_ _02896_ _02827_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08417_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\] _01965_ VGND VGND VPWR
+ VPWR _01966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09397_ _02835_ _02836_ _02772_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08348_ _01891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _01906_ _01907_ _01908_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08279_ _01850_ _01851_ _01748_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10310_ _03625_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _03637_ _03638_ _03633_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11290_ _04491_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10241_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03572_ _03584_
+ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10172_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03523_ VGND
+ VGND VPWR VPWR _03525_ sky130_fd_sc_hd__or2_1
X_14980_ clknet_leaf_95_i_clk _00525_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_13931_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06777_ VGND
+ VGND VPWR VPWR _06778_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13862_ _06715_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12813_ _05809_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__and2_1
X_13793_ _06556_ _06656_ _06657_ _06459_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _05525_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__and2_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12675_ _05670_ _05691_ _05692_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__o31ai_2
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14414_ _07191_ _07192_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__and2_1
X_11626_ _04770_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15394_ clknet_leaf_30_i_clk _00939_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14345_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] VGND VGND VPWR VPWR
+ _07133_ sky130_fd_sc_hd__nor3_1
X_11557_ _04731_ _04729_ _04730_ _04396_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10508_ _03626_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03812_
+ _03813_ _03814_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__o221a_1
X_11488_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__or2_1
X_14276_ _07072_ _07073_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13227_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06136_ VGND
+ VGND VPWR VPWR _06175_ sky130_fd_sc_hd__nor2_1
X_10439_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _03752_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _06112_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__or2b_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _05132_ _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13089_ _06028_ _06050_ net113 _06052_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__a31oi_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07650_ r_i_alpha1\[16\] _01325_ _01258_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__mux2_1
X_07581_ _01259_ _01262_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09320_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__buf_2
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09251_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _02695_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__nor3_1
XFILLER_0_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08202_ _01465_ _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09182_ _02630_ _02632_ _02644_ _02648_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__a31o_2
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08133_ _01691_ _01697_ _01709_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08064_ _01512_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08966_ _02445_ _02448_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nor2_1
X_07917_ _01526_ _01527_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[13\]
+ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__o21a_1
X_08897_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _02376_
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__a211o_1
X_07848_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[3\]
+ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07779_ _01419_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09518_ _02942_ _02933_ _02943_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__a21o_1
X_10790_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _04056_
+ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__nor2_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09449_ _02866_ _02868_ _02876_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a21boi_1
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12460_ _05507_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11411_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12391_ _05139_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _05455_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11342_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] VGND VGND VPWR
+ VPWR _04540_ sky130_fd_sc_hd__inv_2
X_14130_ _06907_ net348 VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11273_ _04477_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
X_14061_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06845_ VGND
+ VGND VPWR VPWR _06893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13012_ _05984_ _05985_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__nand2_2
X_10224_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__clkbuf_4
X_10155_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03508_ VGND
+ VGND VPWR VPWR _03509_ sky130_fd_sc_hd__and2_1
X_14963_ clknet_leaf_95_i_clk _00508_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold6 _00595_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nor2_1
X_13914_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _06716_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__o21a_1
X_14894_ clknet_leaf_109_i_clk _00439_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13845_ _06695_ _06699_ _06694_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13776_ _06642_ _06643_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__o21a_1
X_10988_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _04233_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12727_ _05740_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12658_ _05668_ _05676_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11609_ _04771_ net274 VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15377_ clknet_leaf_29_i_clk _00922_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12589_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05618_ VGND
+ VGND VPWR VPWR _05620_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14328_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _07117_ VGND
+ VGND VPWR VPWR _07118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap114 _05015_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xhold406 _00611_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] VGND VGND VPWR
+ VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR
+ VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold439 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR
+ VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ _07057_ _07058_ _07059_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _02321_ net364 _01945_ _02328_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__o211a_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\] _02264_ _02262_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\]
+ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__a22o_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07702_ _01365_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
X_08682_ _02022_ net574 _02205_ _02206_ _02055_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07633_ diff2\[17\] diff1\[13\] VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07564_ _01257_ diff2\[17\] diff1\[17\] VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09303_ _02754_ net305 _02749_ _02756_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07495_ _01022_ _01138_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09234_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02696_ VGND
+ VGND VPWR VPWR _02697_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09165_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _02634_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08116_ _01708_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__inv_2
X_09096_ _02572_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08047_ _01610_ _01626_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09998_ _03359_ _03364_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__a21oi_1
X_08949_ _01981_ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__and2_1
X_11960_ _05062_ _05065_ _05074_ _05075_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__o31a_1
X_10911_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04150_ _04034_
+ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__o211a_1
X_11891_ _05018_ _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__or2_1
X_13630_ _06516_ _06519_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__nand2_1
X_10842_ _04101_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _04102_ sky130_fd_sc_hd__or2b_1
XFILLER_0_156_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13561_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _06460_ VGND
+ VGND VPWR VPWR _06461_ sky130_fd_sc_hd__and2_1
X_10773_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _04028_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__or3_1
X_15300_ clknet_leaf_19_i_clk _00845_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12512_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _05552_
+ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13492_ _06396_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15231_ clknet_leaf_14_i_clk _00776_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12443_ _05488_ net153 _05495_ _05496_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15162_ clknet_leaf_111_i_clk net238 VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12374_ _05431_ _05434_ _05432_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14113_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _06929_
+ _06934_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__o21ai_1
X_11325_ _04503_ _04524_ _04513_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15093_ clknet_leaf_99_i_clk _00638_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11256_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04460_ VGND
+ VGND VPWR VPWR _04462_ sky130_fd_sc_hd__nand2_1
X_14044_ _06876_ _06877_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10207_ _03517_ _03518_ _03555_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__a21o_1
X_11187_ _04061_ _04398_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nand2_1
X_10138_ _03389_ _03492_ _03493_ _03292_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__o211a_1
X_14946_ clknet_leaf_108_i_clk _00491_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10069_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03410_ VGND
+ VGND VPWR VPWR _03432_ sky130_fd_sc_hd__nand2_1
X_14877_ clknet_leaf_110_i_clk net217 VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13828_ _06688_ _06689_ _06584_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13759_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06628_
+ _06569_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07280_ _01026_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15429_ clknet_leaf_8_i_clk _00974_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold203 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] VGND VGND
+ VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold225 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 r_i_alpha1\[6\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold247 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 net60 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _03296_ VGND
+ VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nand2_1
Xhold269 r_i_alpha1\[15\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _02851_ _03238_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a21bo_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _02315_
+ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _03182_ sky130_fd_sc_hd__inv_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _02234_ _02228_ _02246_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__and3_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\]
+ _02170_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\] _01298_ _01282_ VGND
+ VGND VPWR VPWR _01299_ sky130_fd_sc_hd__mux2_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08596_ _02128_ _02120_ _02121_ _01865_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07547_ net430 net293 _01012_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07478_ _01016_ net302 _01201_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09217_ _02677_ _02680_ _02676_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09148_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02608_ _02342_
+ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09079_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _02555_ _02556_
+ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__nand3_1
X_11110_ _04048_ _04343_ _04344_ _04063_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12090_ _04829_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05177_ _05187_
+ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__o41a_1
X_11041_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _04251_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__or3_1
X_14800_ clknet_leaf_71_i_clk _00345_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12992_ _05848_ net480 VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__or2_1
X_14731_ clknet_leaf_72_i_clk _00276_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_11943_ _04770_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND
+ VGND VPWR VPWR _05068_ sky130_fd_sc_hd__or2_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14662_ clknet_leaf_49_i_clk _00207_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11874_ _04557_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13613_ _06501_ _06507_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10825_ _04085_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14593_ clknet_leaf_49_i_clk _00138_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13544_ _06437_ _06438_ _06436_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__a21o_1
X_10756_ _04023_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _04026_ _04027_ _03814_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13475_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ _06351_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10687_ _03606_ _03974_ _03975_ _03780_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__o211a_1
X_15214_ clknet_leaf_124_i_clk _00759_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12426_ _01529_ _02310_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15145_ clknet_leaf_125_i_clk _00690_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12357_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _05424_ VGND
+ VGND VPWR VPWR _05425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11308_ _04509_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
X_15076_ clknet_leaf_119_i_clk _00621_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12288_ _05290_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__and2_1
X_14027_ _06861_ _06862_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__and2_1
X_11239_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR _04447_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14929_ clknet_leaf_78_i_clk _00474_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08450_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[4\] _01994_ VGND VGND VPWR
+ VPWR _01996_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07401_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _01129_ VGND
+ VGND VPWR VPWR _01138_ sky130_fd_sc_hd__xnor2_1
X_08381_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] _01935_ _01870_
+ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07332_ _01046_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07263_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09002_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02485_ VGND
+ VGND VPWR VPWR _02487_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09904_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _03283_ sky130_fd_sc_hd__inv_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _03184_ _03224_ _03225_ _03058_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__o211a_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _02761_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] VGND
+ VGND VPWR VPWR _03168_ sky130_fd_sc_hd__and2_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _01869_ _02235_ _02236_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09697_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR
+ VPWR _03105_ sky130_fd_sc_hd__inv_2
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _02175_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__inv_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\] _02113_ VGND VGND VPWR
+ VPWR _02114_ sky130_fd_sc_hd__xor2_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ _03650_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__nand2_1
X_11590_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _04758_
+ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10541_ _03828_ _03833_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ _03619_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__clkbuf_4
X_10472_ _03741_ _03742_ _03766_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12211_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _05279_ VGND
+ VGND VPWR VPWR _05295_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13191_ _06141_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ _04850_ _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__and2_1
X_12073_ _05171_ _05173_ _05164_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__mux2_1
X_11024_ _04264_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__nor2_1
X_12975_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05951_ VGND
+ VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14714_ clknet_leaf_53_i_clk _00259_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11926_ _05049_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__and2_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ clknet_leaf_58_i_clk _00190_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _04769_ net312 _04979_ _04988_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10808_ _04048_ _04070_ _04071_ _04063_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14576_ clknet_leaf_41_i_clk _00121_ VGND VGND VPWR VPWR diff1\[1\] sky130_fd_sc_hd__dfxtp_1
X_11788_ _04765_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] VGND
+ VGND VPWR VPWR _04929_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13527_ _06210_ net299 _06203_ _06430_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10739_ _04011_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _04003_ _04013_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13458_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _06370_
+ _06371_ _06285_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12409_ _05463_ _05465_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__a21oi_1
Xoutput105 net105 VGND VGND VPWR VPWR out_sintheta[3] sky130_fd_sc_hd__clkbuf_4
X_13389_ _06307_ _06309_ _06199_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15128_ clknet_leaf_115_i_clk _00673_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15059_ clknet_leaf_112_i_clk _00604_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_07950_ _01539_ net555 _01553_ _01555_ _01513_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__o221a_1
X_07881_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[6\] _01487_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[7\]
+ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__o21ai_1
X_09620_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _03035_ sky130_fd_sc_hd__inv_2
X_09551_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _02973_ VGND
+ VGND VPWR VPWR _02974_ sky130_fd_sc_hd__xor2_2
XFILLER_0_144_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08502_ _02039_ _02042_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__nand2_1
X_09482_ _02911_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08433_ _01980_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08364_ _01550_ _01918_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07315_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _01048_ VGND
+ VGND VPWR VPWR _01061_ sky130_fd_sc_hd__xnor2_1
X_08295_ _01864_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_4
X_07246_ _01002_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09818_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _03204_
+ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nand2_1
X_09749_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03152_ VGND
+ VGND VPWR VPWR _03153_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _05768_ _05771_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__o21a_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _04855_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__nor2_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _05703_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__xor2_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _07156_ VGND
+ VGND VPWR VPWR _07207_ sky130_fd_sc_hd__or2_1
X_11642_ _04798_ _04796_ _04797_ _04755_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14361_ _07143_ _07139_ _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11573_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04746_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 in_alpha[7] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_0_24_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13312_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _06244_
+ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__xnor2_1
X_10524_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__and2_1
Xinput29 in_x[17] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
XFILLER_0_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14292_ _07059_ _07086_ _07087_ _06996_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13243_ _06161_ _06187_ _06188_ _06162_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__a211o_1
X_10455_ _03752_ _03754_ _03747_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13174_ _05845_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nand2_1
X_10386_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _03702_ VGND
+ VGND VPWR VPWR _03704_ sky130_fd_sc_hd__nor2_1
X_12125_ _05215_ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12056_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05148_
+ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__nand2_1
X_11007_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR _04250_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12958_ _05848_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _05937_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11909_ _05033_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12889_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05872_
+ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__o21ai_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14628_ clknet_leaf_58_i_clk _00173_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14559_ clknet_leaf_39_i_clk _00105_ VGND VGND VPWR VPWR diff2\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08080_ _01669_ _01675_ _01470_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08982_ _01981_ _02468_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__and2_1
X_07933_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[15\] _01540_ _01529_
+ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_112_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07864_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[4\]
+ _01469_ _01482_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__o31a_1
X_09603_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _03019_ VGND
+ VGND VPWR VPWR _03020_ sky130_fd_sc_hd__xnor2_1
X_07795_ _01430_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
X_09534_ _02956_ _02952_ _02950_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09465_ _02885_ _02888_ _02894_ _02751_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08416_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[2\] _01964_ VGND VGND VPWR
+ VPWR _01965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09396_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _02830_
+ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08347_ _01512_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08278_ _01718_ net44 _01735_ _01736_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__o31a_1
XFILLER_0_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07229_ _00992_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10240_ _03582_ _03586_ _02132_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10171_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03523_ VGND
+ VGND VPWR VPWR _03524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13930_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__and2b_1
X_13861_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _06716_ _06717_
+ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__a21bo_1
X_12812_ _05806_ _05812_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13792_ _06557_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _06657_ sky130_fd_sc_hd__or2_1
X_12743_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ _05734_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__or3_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_91_i_clk clknet_4_5_0_i_clk VGND VGND VPWR VPWR clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12674_ _05693_ _05694_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__and2_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _07156_ VGND
+ VGND VPWR VPWR _07192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11625_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _04784_
+ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15393_ clknet_leaf_30_i_clk _00938_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14344_ _07122_ _07132_ _01552_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__o21a_1
X_11556_ _04729_ _04730_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10507_ _02308_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14275_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _07042_ _07068_
+ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11487_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR _04669_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13226_ _06163_ _06173_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__and2_1
X_10438_ _03623_ _03750_ _03751_ _03515_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13157_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ _06094_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND
+ VPWR VPWR _06113_ sky130_fd_sc_hd__or4b_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10369_ _03685_ _03687_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__a21oi_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _05203_ sky130_fd_sc_hd__buf_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06010_ VGND
+ VGND VPWR VPWR _06052_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12039_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07580_ _01268_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09250_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND VGND VPWR
+ VPWR _02711_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08201_ _01582_ _01786_ _01329_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09181_ _02621_ _02630_ _02626_ _02644_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__a41o_1
XFILLER_0_145_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08132_ _01709_ _01710_ _01723_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08063_ _01556_ _01659_ _01480_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08965_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02452_ VGND
+ VGND VPWR VPWR _02453_ sky130_fd_sc_hd__xnor2_2
X_07916_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\] _01521_ VGND VGND
+ VPWR VPWR _01527_ sky130_fd_sc_hd__and2b_1
X_08896_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _02383_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__and3_1
X_07847_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[3\]
+ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__nand2_1
X_07778_ _01418_ net404 _01344_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09517_ _02942_ _02933_ _02921_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _02880_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__clkbuf_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _02757_ net623 _02820_ _02821_ _02689_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11410_ _04431_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _04599_
+ _04600_ _04539_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__o221a_1
X_12390_ _05450_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11341_ _04431_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _04536_
+ _04537_ _04539_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14060_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06845_ VGND
+ VGND VPWR VPWR _06892_ sky130_fd_sc_hd__or2_1
X_11272_ _04468_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__and2_1
X_13011_ _05614_ _05983_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__nand2_1
X_10223_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03570_ _03207_
+ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10154_ _03398_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14962_ clknet_leaf_95_i_clk _00507_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold7 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__and2_1
X_13913_ _06717_ _06737_ _06755_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__or4_1
X_14893_ clknet_leaf_78_i_clk _00438_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13844_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _06684_ VGND
+ VGND VPWR VPWR _06703_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13775_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06637_
+ _06587_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__a21oi_1
X_10987_ _04226_ _04224_ _04230_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__or3b_1
X_12726_ _05732_ _05739_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15445_ clknet_leaf_28_i_clk _00990_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12657_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _05648_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11608_ _04770_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15376_ clknet_leaf_29_i_clk _00921_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05618_ VGND
+ VGND VPWR VPWR _05619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14327_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _07116_ VGND
+ VGND VPWR VPWR _07117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11539_ _04695_ _04698_ _04707_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold407 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold418 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14258_ _06903_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__clkbuf_4
Xhold429 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND VPWR VPWR
+ net546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13209_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06112_ VGND
+ VGND VPWR VPWR _06159_ sky130_fd_sc_hd__nand2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _06905_ _06997_ _06998_ _06996_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__o211a_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _02267_
+ _02268_ _02055_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__o221a_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ net345 _01364_ _01358_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__mux2_1
X_08681_ _02199_ _02195_ _02204_ _01924_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__a31o_1
X_07632_ _01311_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07563_ diff3\[17\] VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09302_ _02755_ net356 VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07494_ _01015_ net505 _01212_ _01213_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09233_ _02343_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09164_ _02621_ _02626_ _02632_ _02630_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08115_ _01706_ _01707_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09095_ _02497_ _02571_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08046_ _01643_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09997_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _03366_ VGND
+ VGND VPWR VPWR _03367_ sky130_fd_sc_hd__xnor2_2
X_08948_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02437_ _02319_
+ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__mux2_1
X_08879_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _02378_
+ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__xnor2_1
X_10910_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR _04164_ sky130_fd_sc_hd__inv_2
X_11890_ _05014_ _05017_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10841_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04100_ VGND
+ VGND VPWR VPWR _04101_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06410_ VGND
+ VGND VPWR VPWR _06460_ sky130_fd_sc_hd__nor2_1
X_10772_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04018_ VGND VGND
+ VPWR VPWR _04041_ sky130_fd_sc_hd__and4_1
X_12511_ _05203_ _05549_ _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13491_ _06397_ _06398_ _06399_ _06388_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15230_ clknet_leaf_15_i_clk _00775_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12442_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] _05492_
+ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15161_ clknet_leaf_55_i_clk _00706_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
X_12373_ _05437_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14112_ _06646_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__inv_2
X_11324_ _04511_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _04524_ sky130_fd_sc_hd__or2b_1
X_15092_ clknet_leaf_120_i_clk _00637_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14043_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06845_ VGND
+ VGND VPWR VPWR _06877_ sky130_fd_sc_hd__nand2_1
X_11255_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04460_ VGND
+ VGND VPWR VPWR _04461_ sky130_fd_sc_hd__or2_1
X_10206_ _03526_ _03531_ _03539_ _03548_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__or4_1
X_11186_ _04390_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _04401_ _04402_ _04360_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__o221a_1
X_10137_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND
+ VGND VPWR VPWR _03493_ sky130_fd_sc_hd__or2_1
X_14945_ clknet_leaf_109_i_clk _00490_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10068_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03410_ VGND
+ VGND VPWR VPWR _03431_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14876_ clknet_leaf_78_i_clk _00421_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13827_ _06671_ _06679_ _06687_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13758_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06628_
+ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12709_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _05723_ VGND
+ VGND VPWR VPWR _05725_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13689_ _06565_ net524 _06568_ _06570_ _06526_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15428_ clknet_leaf_9_i_clk _00973_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15359_ clknet_leaf_19_i_clk _00904_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold204 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold215 r_i_alpha1\[5\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _00657_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 r_i_alpha1\[13\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09920_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _03296_ VGND
+ VGND VPWR VPWR _03297_ sky130_fd_sc_hd__or2_1
Xhold248 r_i_alpha1\[4\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold259 r_i_alpha1\[16\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09851_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _03228_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _03239_ sky130_fd_sc_hd__a31o_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _02315_ sky130_fd_sc_hd__clkbuf_4
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _03181_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__clkbuf_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _02213_ _02222_ _02234_ _02246_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__and4bb_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _02173_ _02183_ _02184_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07615_ r_i_alpha1\[9\] _01297_ _01276_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__mux2_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08595_ _02120_ _02121_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07546_ _01245_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07477_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _01159_ _01199_
+ _01200_ _01030_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09216_ _02676_ _02677_ _02680_ _02313_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09147_ _02329_ net473 _02381_ _02617_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09078_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _02553_ VGND
+ VGND VPWR VPWR _02556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08029_ net35 net53 VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11040_ _04279_ _04274_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12991_ _05960_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11942_ _05065_ _05066_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__nor2_1
X_14730_ clknet_leaf_73_i_clk _00275_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ clknet_leaf_58_i_clk _00206_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04794_ VGND VGND VPWR
+ VPWR _05003_ sky130_fd_sc_hd__o31a_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13612_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06506_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__mux2_1
X_10824_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04084_ VGND
+ VGND VPWR VPWR _04086_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14592_ clknet_leaf_38_i_clk _00137_ VGND VGND VPWR VPWR diff3\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13543_ _06443_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__or2b_1
XFILLER_0_149_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10755_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04025_
+ _04012_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13474_ _06365_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__nand2_1
X_10686_ _03608_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] VGND
+ VGND VPWR VPWR _03975_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15213_ clknet_leaf_2_i_clk _00758_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_35_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12425_ net536 _05140_ _05482_ _05483_ _05391_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__o221a_1
XFILLER_0_51_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15144_ clknet_leaf_125_i_clk _00689_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12356_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _05420_ _05423_
+ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _04468_ _04508_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15075_ clknet_leaf_100_i_clk _00620_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12287_ _05139_ _05357_ _05358_ _05360_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14026_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06837_ VGND
+ VGND VPWR VPWR _06862_ sky130_fd_sc_hd__nand2_1
X_11238_ _04442_ _04443_ _04446_ _04063_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11169_ _04379_ net274 VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14928_ clknet_leaf_81_i_clk _00473_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14859_ clknet_leaf_86_i_clk _00404_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07400_ _01095_ net197 _01136_ _01137_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\] _01935_ VGND VGND
+ VPWR VPWR _01936_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07331_ _01016_ net284 _01074_ _01075_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07262_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _01012_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09001_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02485_ VGND
+ VGND VPWR VPWR _02486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09903_ _03189_ _03280_ _03017_ _03282_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09834_ net124 _03190_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__or2_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _02755_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03166_
+ _03167_ _03013_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__o221a_1
X_08716_ _01868_ _02237_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__nor2_1
X_09696_ _02748_ _03103_ _03104_ _03058_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__o211a_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _02173_ _02174_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__or2_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08578_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[16\] _02112_ VGND VGND VPWR
+ VPWR _02113_ sky130_fd_sc_hd__xnor2_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07529_ net434 net215 _01234_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10540_ _03832_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _03842_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10471_ _03765_ _03776_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12210_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _05279_ VGND
+ VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13190_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06142_ _06138_
+ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12141_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _05231_ _01249_
+ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12072_ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__inv_2
X_11023_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _04263_ VGND
+ VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nor2_1
X_12974_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05950_ VGND
+ VGND VPWR VPWR _05951_ sky130_fd_sc_hd__xnor2_1
X_14713_ clknet_leaf_50_i_clk net470 VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11925_ _05050_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11856_ _04986_ _04987_ _04786_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__o21ai_1
X_14644_ clknet_leaf_59_i_clk _00189_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _04010_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _04071_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14575_ clknet_leaf_41_i_clk _00120_ VGND VGND VPWR VPWR diff1\[0\] sky130_fd_sc_hd__dfxtp_1
X_11787_ _04925_ _04927_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10738_ _04012_ net258 VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__nand2_1
X_13526_ _06232_ _06429_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13457_ _06362_ _06365_ _06369_ _06205_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__o31ai_1
X_10669_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03944_ VGND
+ VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12408_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05423_ VGND
+ VGND VPWR VPWR _05469_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13388_ _06296_ _06300_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__o21a_1
Xoutput106 net106 VGND VGND VPWR VPWR out_sintheta[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15127_ clknet_leaf_116_i_clk _00672_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12339_ _05403_ _05406_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__and2_1
X_15058_ clknet_leaf_112_i_clk _00603_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14009_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _06848_ sky130_fd_sc_hd__or2_1
X_07880_ _01463_ net546 _01460_ _01496_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__o211a_1
X_09550_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _02964_ _02772_
+ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__o21a_1
X_08501_ _02039_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__or2_1
X_09481_ _02497_ _02910_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08432_ _01978_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08363_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[9\] _01914_ _01916_
+ _01550_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__a2bb2o_1
X_07314_ _01044_ net171 _01060_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08294_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_out VGND VGND VPWR VPWR _01864_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07245_ net338 net5 _01000_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09817_ net266 _03189_ _03017_ _03210_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03149_ _03151_
+ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__a21oi_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03088_ VGND
+ VGND VPWR VPWR _03089_ sky130_fd_sc_hd__xor2_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _04844_ _04846_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__nand2_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12690_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _05707_ VGND
+ VGND VPWR VPWR _05708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _04796_ _04797_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a21oi_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14360_ _07145_ _07146_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11572_ _04742_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13311_ _06241_ _06243_ _06235_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__mux2_1
X_10523_ _03626_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03826_
+ _03827_ _03814_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__o221a_1
Xinput19 in_alpha[8] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
X_14291_ _06909_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND
+ VGND VPWR VPWR _07087_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13242_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _06142_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__o41a_1
X_10454_ _03749_ _03755_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13173_ _06115_ _06123_ _06126_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__o21ai_1
X_10385_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _03702_ VGND
+ VGND VPWR VPWR _03703_ sky130_fd_sc_hd__and2_1
X_12124_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05214_ VGND
+ VGND VPWR VPWR _05216_ sky130_fd_sc_hd__nand2_1
X_12055_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _05145_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__or3_1
X_11006_ _04249_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12957_ _05931_ _05935_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11908_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05034_ VGND
+ VGND VPWR VPWR _05035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14627_ clknet_leaf_59_i_clk _00172_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_11839_ _04850_ _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14558_ clknet_leaf_37_i_clk _00104_ VGND VGND VPWR VPWR diff1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13509_ _06414_ _06415_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14489_ clknet_leaf_5_i_clk _00035_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08981_ _02313_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02466_
+ _02467_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07932_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[15\] _01540_ VGND VGND
+ VPWR VPWR _01541_ sky130_fd_sc_hd__and2_1
X_07863_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[17\] _01476_ VGND VGND
+ VPWR VPWR _01482_ sky130_fd_sc_hd__nand2_1
X_09602_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _03018_ VGND
+ VGND VPWR VPWR _03019_ sky130_fd_sc_hd__xnor2_1
X_07794_ net390 _01429_ _01411_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__mux2_1
X_09533_ _02956_ _02952_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09464_ _02885_ _02888_ _02894_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08415_ _01549_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR _01964_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09395_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _02829_
+ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08346_ _01905_ _01903_ _01904_ _01870_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_148_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08277_ _01758_ _01830_ _01839_ _01756_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07228_ net2 VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10170_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03522_ VGND
+ VGND VPWR VPWR _03523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13860_ _06710_ _06711_ _06708_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__a21bo_1
X_12811_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _05789_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__o21a_1
X_13791_ _06651_ _06655_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _05755_ sky130_fd_sc_hd__inv_2
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05648_ VGND
+ VGND VPWR VPWR _05694_ sky130_fd_sc_hd__nand2_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _04445_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _04775_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__o31a_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _07144_ VGND
+ VGND VPWR VPWR _07191_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15392_ clknet_leaf_27_i_clk net246 VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11555_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04723_ VGND
+ VGND VPWR VPWR _04731_ sky130_fd_sc_hd__xnor2_1
X_14343_ _07130_ _07131_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10506_ _03805_ _03808_ _03811_ _03631_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__a31o_1
X_14274_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _07041_ VGND
+ VGND VPWR VPWR _07072_ sky130_fd_sc_hd__xnor2_1
X_11486_ _04431_ net406 _04667_ _04668_ _04539_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__o221a_1
X_13225_ _06160_ _06168_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__and2_1
X_10437_ _03621_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _03751_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13156_ _06111_ _05566_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__mux2_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _03685_ _03687_ _03642_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__o21ai_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05198_
+ _05197_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a21oi_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _06010_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__o41ai_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__or2_1
X_12038_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13989_ _06820_ _06823_ _06821_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08200_ _01579_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09180_ _02638_ _02641_ _02643_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08131_ net25 net43 VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08062_ _01653_ _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08964_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _02451_ VGND
+ VGND VPWR VPWR _02452_ sky130_fd_sc_hd__xor2_2
X_07915_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\] _01523_ VGND VGND
+ VPWR VPWR _01526_ sky130_fd_sc_hd__and2_1
X_08895_ net481 VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07846_ _01464_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07777_ _01334_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__inv_2
X_09516_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND VPWR
+ VPWR _02942_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09447_ _02497_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__and2_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09378_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _02818_
+ _02819_ _02761_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08329_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND VPWR VPWR _01892_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11340_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11271_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04475_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13010_ _05614_ _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__or2_1
X_10222_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03569_ VGND
+ VGND VPWR VPWR _03570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10153_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03206_ _03495_
+ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14961_ clknet_leaf_90_i_clk _00506_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_10084_ _03389_ _03444_ _03445_ _03292_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__o211a_1
Xhold8 _00430_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
X_13912_ _06736_ _06743_ _06748_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__or3b_1
X_14892_ clknet_leaf_109_i_clk _00437_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13843_ _06702_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10986_ _04226_ _04224_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13774_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _06632_ _06587_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12725_ _05732_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15444_ clknet_leaf_27_i_clk _00989_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12656_ _05487_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] VGND
+ VGND VPWR VPWR _05679_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_111_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_111_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11607_ _04757_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__buf_2
X_12587_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05617_ VGND
+ VGND VPWR VPWR _05618_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15375_ clknet_leaf_29_i_clk _00920_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14326_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__and2b_1
X_11538_ _04678_ _04679_ _04715_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND VPWR
+ VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _04631_ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__or2_1
X_14257_ _07056_ _07054_ _07055_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13208_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06136_ VGND
+ VGND VPWR VPWR _06158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14188_ _06907_ net412 VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__or2_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _06096_ VGND
+ VGND VPWR VPWR _06097_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ net7 _01361_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__xor2_1
X_08680_ _02199_ _02195_ _02204_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__a21oi_1
X_07631_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\] _01310_ _01282_
+ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07562_ _01256_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09301_ _02750_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__clkbuf_4
X_07493_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _01045_ _01013_
+ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09232_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _02671_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09163_ _02599_ _02603_ _02614_ _02622_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08114_ net25 net43 VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09094_ _02319_ _02568_ _02569_ _02570_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08045_ _01612_ _01627_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_i_clk clknet_4_5_0_i_clk VGND VGND VPWR VPWR clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09996_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03365_ VGND
+ VGND VPWR VPWR _03366_ sky130_fd_sc_hd__xor2_2
X_08947_ _02435_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08878_ _01959_ _02376_ _02377_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__o21ai_1
X_07829_ _01251_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_4
X_10840_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04093_ _04033_
+ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10771_ _04023_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04039_ _04040_ _03814_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__o221a_1
X_12510_ _05203_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nand2_1
X_13490_ _06383_ _06393_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12441_ _03619_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12372_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05430_ VGND
+ VGND VPWR VPWR _05438_ sky130_fd_sc_hd__nand2_1
X_15160_ clknet_leaf_122_i_clk _00705_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11323_ _04521_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__and2_1
X_14111_ _06928_ net316 _06932_ _06933_ _06922_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15091_ clknet_leaf_99_i_clk _00636_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11254_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04459_ VGND
+ VGND VPWR VPWR _04460_ sky130_fd_sc_hd__xnor2_1
X_14042_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06845_ VGND
+ VGND VPWR VPWR _06876_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10205_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03547_ _03553_
+ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11185_ _04395_ _04400_ _04376_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10136_ _03490_ _03491_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14944_ clknet_leaf_107_i_clk net259 VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10067_ _03389_ _03429_ _03430_ _03292_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14875_ clknet_leaf_75_i_clk _00420_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13826_ _06671_ _06679_ _06687_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13757_ _06626_ _06627_ _06587_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__mux2_1
X_10969_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12708_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _05723_ VGND
+ VGND VPWR VPWR _05724_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13688_ _06293_ _06566_ _06567_ _06569_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__a31o_1
X_15427_ clknet_leaf_26_i_clk _00972_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12639_ _05655_ _05658_ _05663_ _05487_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ clknet_leaf_19_i_clk _00903_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14309_ _07057_ _07079_ _07096_ _07101_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__or4_1
Xhold205 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold216 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ clknet_leaf_17_i_clk _00834_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold227 r_i_alpha1\[10\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold249 net61 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _03233_
+ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__or2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__buf_4
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _02751_ _02310_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__and2_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\] _02251_ VGND VGND VPWR
+ VPWR _02252_ sky130_fd_sc_hd__xor2_2
X_08663_ _02177_ _02185_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07614_ diff2\[9\] _01270_ _01272_ diff3\[9\] _01296_ VGND VGND VPWR VPWR _01297_
+ sky130_fd_sc_hd__a221o_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _02126_ _02127_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__or2_1
X_07545_ net415 net278 _01012_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07476_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _01122_ _01101_
+ _01047_ _01072_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09215_ _02649_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09146_ _02615_ _02616_ _02320_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09077_ _02554_ _02344_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__mux2_2
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08028_ _01625_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09979_ _03184_ _03349_ _03350_ _03292_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__o211a_1
X_12990_ _05964_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11941_ _05064_ _05056_ _05058_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__and3_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ clknet_leaf_58_i_clk _00205_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _05002_ sky130_fd_sc_hd__inv_2
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06504_ _06505_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10823_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _04084_ VGND
+ VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nand2_1
X_14591_ clknet_leaf_37_i_clk _00136_ VGND VGND VPWR VPWR diff3\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13542_ _06080_ _06442_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__nand2_1
X_10754_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _04025_
+ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10685_ _03972_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__xnor2_1
X_13473_ _06369_ _06375_ _06379_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__nor3_1
XFILLER_0_125_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15212_ clknet_leaf_2_i_clk _00757_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_12424_ _05473_ _05477_ _05481_ _05222_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15143_ clknet_leaf_125_i_clk _00688_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12355_ _05422_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11306_ _04375_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04506_
+ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__a22o_1
X_15074_ clknet_leaf_119_i_clk _00619_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_12286_ _01249_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11237_ _04444_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__or2_1
X_14025_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _06837_ VGND
+ VGND VPWR VPWR _06861_ sky130_fd_sc_hd__or2_1
X_11168_ _04377_ net276 _04387_ _04388_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10119_ _03468_ _03471_ _03467_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__a21oi_2
X_11099_ _04328_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__inv_2
X_14927_ clknet_leaf_81_i_clk _00472_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14858_ clknet_leaf_85_i_clk _00403_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13809_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _06670_ VGND
+ VGND VPWR VPWR _06672_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14789_ clknet_leaf_66_i_clk _00334_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_07330_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _01029_ _01030_
+ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07261_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ _01010_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09000_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _02484_ VGND
+ VGND VPWR VPWR _02485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09902_ _03277_ _03281_ _03191_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _03223_
+ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__xnor2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _03162_ _03159_ _03165_ _02751_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__o31ai_1
X_08715_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] VGND VGND VPWR
+ VPWR _02237_ sky130_fd_sc_hd__inv_2
X_09695_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _03104_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _02169_ _02172_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__and2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _01882_ _02111_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__and2_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07528_ _01236_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07459_ _01022_ _01061_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10470_ _03623_ _03778_ _03779_ _03780_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09129_ _02599_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12140_ _05229_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12071_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _05158_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__or3_1
X_11022_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _04263_ VGND
+ VGND VPWR VPWR _04264_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12973_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05877_ VGND VGND
+ VPWR VPWR _05950_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14712_ clknet_leaf_50_i_clk _00257_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11924_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _05048_ VGND
+ VGND VPWR VPWR _05050_ sky130_fd_sc_hd__nor2_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ clknet_leaf_59_i_clk _00188_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _04980_ _04985_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__and2_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ _04065_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14574_ clknet_leaf_39_i_clk net2 VGND VGND VPWR VPWR diff_valid sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11786_ _04907_ _04910_ _04918_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13525_ _06421_ _06428_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__xnor2_1
X_10737_ _04010_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13456_ _06362_ _06365_ _06369_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10668_ _03957_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12407_ _05468_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10599_ _03608_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND
+ VGND VPWR VPWR _03896_ sky130_fd_sc_hd__or2_1
X_13387_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _06299_ VGND
+ VGND VPWR VPWR _06308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR out_sintheta[5] sky130_fd_sc_hd__clkbuf_4
X_15126_ clknet_leaf_116_i_clk _00671_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12338_ _05403_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15057_ clknet_leaf_108_i_clk _00602_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12269_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14008_ _06844_ _06846_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08500_ _01998_ _02005_ _02014_ _02030_ _02041_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__a41o_1
X_09480_ _02746_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _02908_
+ _02909_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08431_ _01251_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08362_ _01891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _01919_ _01920_ _01908_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07313_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _01045_ _01050_
+ _01058_ _01059_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__o221a_1
X_08293_ _01863_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07244_ _01001_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09816_ _03191_ _03209_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__nand2_1
X_09747_ _03150_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR VPWR
+ _03151_ sky130_fd_sc_hd__mux2_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _02771_ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__nand2_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR VPWR
+ _02158_ sky130_fd_sc_hd__inv_2
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] VGND VGND
+ VPWR VPWR _04798_ sky130_fd_sc_hd__inv_2
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11571_ _04730_ _04743_ _04744_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13310_ _06242_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10522_ _03816_ _03821_ _03825_ _03631_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14290_ _07084_ _07085_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13241_ _06177_ _06173_ _06181_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__and3_1
X_10453_ _03763_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13172_ _06115_ _06123_ _06126_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nor3_1
X_10384_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03701_ VGND
+ VGND VPWR VPWR _03702_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12123_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05214_ VGND
+ VGND VPWR VPWR _05215_ sky130_fd_sc_hd__nor2_1
X_12054_ _05153_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _05156_ _05157_ _04965_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__o221a_1
X_11005_ _04248_ _03118_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12956_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _05934_ VGND
+ VGND VPWR VPWR _05935_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11907_ _04952_ net114 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__a21oi_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _05877_ sky130_fd_sc_hd__inv_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ clknet_leaf_59_i_clk _00171_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_11838_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04972_ _04757_
+ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14557_ clknet_leaf_37_i_clk _00103_ VGND VGND VPWR VPWR diff1\[16\] sky130_fd_sc_hd__dfxtp_1
X_11769_ _04910_ _04911_ _04862_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13508_ _06387_ _06413_ _06412_ _06200_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14488_ clknet_leaf_5_i_clk _00034_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13439_ _06350_ _06353_ _06205_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15109_ clknet_leaf_110_i_clk net163 VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_08980_ _02465_ _02457_ _02460_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07931_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[14\] _01532_ _01537_
+ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__o21ai_1
X_07862_ _01467_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[4\] _01479_
+ _01481_ _01475_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__o221a_1
X_09601_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07793_ _01427_ _01428_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09532_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR
+ VPWR _02956_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09463_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02893_ VGND
+ VGND VPWR VPWR _02894_ sky130_fd_sc_hd__xor2_2
XFILLER_0_59_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08414_ _01891_ net465 _01962_ _01963_ _01908_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__o221a_1
X_09394_ _02754_ net547 _02749_ _02834_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__o211a_1
X_08345_ _01903_ _01904_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08276_ _01330_ _01755_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07227_ net15 VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12810_ _05632_ _05814_ _05815_ _05675_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13790_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _06654_ VGND
+ VGND VPWR VPWR _06655_ sky130_fd_sc_hd__xnor2_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _05737_ _05746_ _05747_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__o21ai_2
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05648_ VGND
+ VGND VPWR VPWR _05693_ sky130_fd_sc_hd__or2_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _06911_ net549 _07189_ _07190_ _01456_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__o221a_1
X_11623_ _04445_ _04778_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__nand2_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ clknet_leaf_23_i_clk _00936_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14342_ _07123_ _07120_ _07129_ _06926_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__a31o_1
X_11554_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _04723_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10505_ _03805_ _03808_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14273_ _07071_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
X_11485_ _04660_ _04657_ _04666_ _04391_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_107_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13224_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _06142_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__o21a_1
X_10436_ _03743_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13155_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ _06094_ _05877_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__o31a_1
X_10367_ _03672_ _03676_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__o21ai_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _05153_ net485 _05200_ _05201_ _05170_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__o221a_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _06027_ _06037_ _06038_ _06044_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__or4_1
X_10298_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nand2_1
X_12037_ _05140_ net342 _05141_ _05143_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13988_ _06827_ _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12939_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05917_
+ _05878_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14609_ clknet_leaf_46_i_clk _00154_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08130_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08061_ _01638_ _01647_ _01637_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08963_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _02442_ _02341_
+ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07914_ _01467_ net559 _01524_ _01525_ _01513_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__o221a_1
X_08894_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _02390_ _02391_ _02309_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__o221a_1
X_07845_ _01463_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\] _01460_
+ _01466_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07776_ _01417_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09515_ _02940_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09446_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02878_ _02750_
+ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__mux2_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09377_ _02818_ _02819_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08328_ _01869_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08259_ _01709_ _01834_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11270_ _04473_ _04474_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10221_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _03536_ VGND VGND
+ VPWR VPWR _03569_ sky130_fd_sc_hd__nor4_2
X_10152_ _03506_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
X_14960_ clknet_leaf_90_i_clk _00505_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10083_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _03445_ sky130_fd_sc_hd__or2_1
Xhold9 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ _06759_ _06760_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__nand2_1
X_14891_ clknet_leaf_78_i_clk _00436_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13842_ _06501_ _06701_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13773_ _06565_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _06640_ _06641_ _06631_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__o221a_1
X_10985_ _04227_ _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__xnor2_1
X_12724_ _05737_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15443_ clknet_leaf_30_i_clk _00988_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_128_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12655_ _05521_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05677_
+ _05678_ _05544_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11606_ _04765_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__clkbuf_4
X_15374_ clknet_leaf_29_i_clk _00919_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12586_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _05598_ _05526_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14325_ _06910_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] _01766_
+ _07115_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11537_ _04676_ _04685_ _04695_ _04707_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__or4_4
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap117 _03700_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_1
Xhold409 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ _07054_ _07055_ _07056_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__o21ai_2
X_11468_ _04635_ _04640_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13207_ _05855_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _06156_
+ _06157_ _05910_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10419_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _03733_ VGND
+ VGND VPWR VPWR _03734_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14187_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _06992_
+ _06991_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__a21oi_1
X_11399_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04565_ VGND
+ VGND VPWR VPWR _04591_ sky130_fd_sc_hd__or2_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06095_ VGND
+ VGND VPWR VPWR _06096_ sky130_fd_sc_hd__xor2_2
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] VGND
+ VGND VPWR VPWR _06036_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07630_ r_i_alpha1\[12\] _01309_ _01276_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__mux2_1
X_07561_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_1
X_09300_ _02751_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07492_ _01076_ _01134_ _01131_ _01080_ _01211_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__a221o_1
X_09231_ _02649_ _02679_ _02690_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09162_ _02615_ _02626_ _02630_ _02621_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08113_ net43 net25 VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__nand2b_1
X_09093_ _02312_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] VGND
+ VGND VPWR VPWR _02570_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08044_ _01638_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09995_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03356_ _03206_
+ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08946_ _02424_ _02427_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08877_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02371_
+ _01959_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__o21ai_1
X_07828_ _01453_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_4
X_07759_ net8 _01400_ net9 VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10770_ _04038_ _04036_ _04037_ _03994_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09429_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND VPWR
+ VPWR _02863_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12440_ _05488_ net149 _05141_ _05494_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12371_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _05430_ VGND
+ VGND VPWR VPWR _05437_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14110_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _06931_
+ _01862_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__o21ai_1
X_11322_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04520_ VGND
+ VGND VPWR VPWR _04522_ sky130_fd_sc_hd__or2_1
X_15090_ clknet_leaf_120_i_clk _00635_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14041_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND VGND
+ VPWR VPWR _06875_ sky130_fd_sc_hd__inv_2
X_11253_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ _04061_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__o21ba_1
X_10204_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03547_ _03549_
+ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11184_ _04395_ _04400_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__nor2_1
X_10135_ _03476_ _03482_ _03480_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__o21a_1
X_14943_ clknet_leaf_109_i_clk _00488_ VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10066_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND
+ VGND VPWR VPWR _03430_ sky130_fd_sc_hd__or2_1
X_14874_ clknet_leaf_79_i_clk _00419_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_13825_ _06685_ _06686_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13756_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _06616_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__or3_1
X_10968_ _04213_ _04214_ _04215_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12707_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05722_ VGND
+ VGND VPWR VPWR _05723_ sky130_fd_sc_hd__xor2_1
Xclkbuf_4_12_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_12_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13687_ _06554_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__clkbuf_4
X_10899_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04152_ VGND
+ VGND VPWR VPWR _04154_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15426_ clknet_leaf_28_i_clk _00971_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12638_ _05655_ _05658_ _05663_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15357_ clknet_leaf_20_i_clk _00902_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12569_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _05600_ VGND
+ VGND VPWR VPWR _05602_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14308_ _07088_ _07090_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15288_ clknet_leaf_14_i_clk _00833_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold206 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold217 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 diff1\[13\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14239_ _07041_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__clkbuf_4
Xhold239 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND
+ VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _02312_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__clkbuf_4
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _02747_ _03179_ _03180_ _03058_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__o211a_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\] _02250_ VGND VGND VPWR
+ VPWR _02251_ sky130_fd_sc_hd__xnor2_2
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _01866_ _02187_ _02188_ _01552_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__o211a_1
X_07613_ _01273_ diff1\[9\] VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[16\] _02125_ VGND VGND VPWR
+ VPWR _02127_ sky130_fd_sc_hd__nor2_1
X_07544_ _01244_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07475_ _01080_ _01096_ _01097_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09214_ _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09145_ _02599_ _02603_ _02614_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nor3_1
XFILLER_0_133_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09076_ _01958_ _02553_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08027_ net36 _01624_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09978_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _03350_ sky130_fd_sc_hd__or2_1
X_08929_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _02416_ VGND
+ VGND VPWR VPWR _02420_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_110_i_clk clknet_4_3_0_i_clk VGND VGND VPWR VPWR clknet_leaf_110_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11940_ _05056_ _05058_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _04990_ _04992_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__or2_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _06495_ _06496_ _06497_ _06490_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_125_i_clk clknet_4_0_0_i_clk VGND VGND VPWR VPWR clknet_leaf_125_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10822_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04083_ VGND
+ VGND VPWR VPWR _04084_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14590_ clknet_leaf_37_i_clk _00135_ VGND VGND VPWR VPWR diff3\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13541_ _06080_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10753_ _03669_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _04015_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__o31a_1
XFILLER_0_95_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13472_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06351_ VGND
+ VGND VPWR VPWR _06383_ sky130_fd_sc_hd__xnor2_1
X_10684_ _03967_ _03968_ _03965_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15211_ clknet_leaf_124_i_clk _00756_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_12423_ _05473_ _05477_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15142_ clknet_leaf_125_i_clk _00687_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12354_ _05421_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR VPWR
+ _05422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11305_ _04505_ _04498_ _04499_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__o31a_1
X_15073_ clknet_leaf_118_i_clk _00618_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12285_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _05359_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14024_ _06563_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _06859_
+ _06860_ _06631_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__o221a_1
X_11236_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _04445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11167_ net161 _04379_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__or2_1
X_10118_ _03475_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
X_11098_ _04319_ _04309_ _04327_ _04328_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14926_ clknet_leaf_82_i_clk _00471_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_10049_ _03394_ _03403_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14857_ clknet_leaf_79_i_clk _00402_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13808_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _06670_ VGND
+ VGND VPWR VPWR _06671_ sky130_fd_sc_hd__nand2_1
X_14788_ clknet_leaf_67_i_clk _00333_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_133_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13739_ _06607_ _06612_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07260_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR _01010_ sky130_fd_sc_hd__buf_2
XFILLER_0_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15409_ clknet_leaf_32_i_clk _00954_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09901_ _03276_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _02851_ _03221_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__o21ai_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _03162_ _03159_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__o21a_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _02234_ _02228_ _02230_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__or3b_1
X_09694_ _03099_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__xnor2_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _02169_ _02172_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\] _02083_ VGND VGND VPWR VPWR
+ _02111_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07527_ net417 net339 _01234_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_i_clk clknet_4_15_0_i_clk VGND VGND VPWR VPWR clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07458_ _01095_ net609 _01185_ _01186_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07389_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09128_ _02156_ _02598_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09059_ _02387_ net644 _02537_ _02538_ _02414_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12070_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05148_ VGND VGND
+ VPWR VPWR _05171_ sky130_fd_sc_hd__and4_1
X_11021_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04262_ VGND
+ VGND VPWR VPWR _04263_ sky130_fd_sc_hd__xor2_1
X_12972_ _05949_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
X_11923_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _05048_ VGND
+ VGND VPWR VPWR _05049_ sky130_fd_sc_hd__nand2_1
X_14711_ clknet_leaf_50_i_clk _00256_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ clknet_leaf_59_i_clk _00187_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _04980_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__nor2_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _04068_ VGND
+ VGND VPWR VPWR _04069_ sky130_fd_sc_hd__xnor2_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14573_ clknet_leaf_36_i_clk _00119_ VGND VGND VPWR VPWR diff2\[17\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11785_ _04917_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13524_ _06426_ _06427_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__nor2_1
X_10736_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13455_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _06351_ VGND
+ VGND VPWR VPWR _06369_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10667_ _03948_ _03950_ _03946_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12406_ _05290_ _05467_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ _06305_ _06306_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__or2b_1
X_10598_ _03893_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15125_ clknet_leaf_116_i_clk _00670_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12337_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05405_ VGND
+ VGND VPWR VPWR _05406_ sky130_fd_sc_hd__xor2_1
Xoutput108 net108 VGND VGND VPWR VPWR out_sintheta[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15056_ clknet_leaf_112_i_clk net275 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12268_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14007_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06845_ _06839_
+ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__a21oi_1
X_11219_ _04390_ net359 _04387_ _04430_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12199_ _05140_ net640 _05141_ _05284_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput90 net90 VGND VGND VPWR VPWR out_costheta[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14909_ clknet_leaf_82_i_clk _00454_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_08430_ _01865_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _01976_
+ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08361_ _01918_ _01915_ _01917_ _01870_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07312_ _01012_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ _01862_ _01253_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07243_ net344 net4 _01000_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09815_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _03208_
+ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09746_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _03149_
+ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _03069_ _03086_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__or2_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _02146_ _02148_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _02082_ _02088_ _02086_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11570_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _04723_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10521_ _03816_ _03821_ _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13240_ _06184_ _06185_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10452_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03762_ VGND
+ VGND VPWR VPWR _03764_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13171_ _06124_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10383_ _03280_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nor2_1
X_12122_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05213_ VGND
+ VGND VPWR VPWR _05214_ sky130_fd_sc_hd__xnor2_1
X_12053_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05155_
+ _01250_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__o21ai_1
X_11004_ _03996_ _04237_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__o21a_1
X_12955_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05933_ VGND
+ VGND VPWR VPWR _05934_ sky130_fd_sc_hd__xnor2_1
X_11906_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _05033_ sky130_fd_sc_hd__inv_2
X_12886_ _05871_ net553 _05875_ _05876_ _05751_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__o221a_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11837_ _04968_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__xnor2_1
X_14625_ clknet_leaf_59_i_clk _00170_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ clknet_leaf_37_i_clk _00102_ VGND VGND VPWR VPWR diff1\[15\] sky130_fd_sc_hd__dfxtp_1
X_11768_ _04909_ _04901_ _04902_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10719_ _03995_ net225 _03620_ _04001_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__o211a_1
X_13507_ _06387_ _06412_ _06413_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__a21oi_1
X_14487_ clknet_leaf_4_i_clk _00033_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ _04754_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04846_
+ _04847_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_43_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13438_ _06350_ _06353_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer1 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND
+ VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13369_ _06292_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15108_ clknet_leaf_111_i_clk _00653_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_15039_ clknet_leaf_96_i_clk _00584_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_07930_ _01464_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07861_ _01471_ _01478_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__a21o_1
X_09600_ _01455_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07792_ net18 net19 _01423_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09531_ _02844_ net521 _02954_ _02955_ _02827_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__o221a_1
X_09462_ _02891_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__xnor2_2
X_08413_ _01961_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[0\] _01866_ VGND
+ VGND VPWR VPWR _01963_ sky130_fd_sc_hd__a21o_1
X_09393_ _02828_ _02832_ _02833_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08344_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND VPWR VPWR
+ _01905_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08275_ _01717_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[15\] _01823_ _01848_
+ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09729_ _03110_ _03124_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12740_ _05732_ _05752_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__or2_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _05648_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__o41a_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _07182_ _07184_ _07188_ _06926_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__a31o_1
X_11622_ _04773_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ _04781_ _04782_ _04539_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ clknet_leaf_23_i_clk _00935_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14341_ _07123_ _07120_ _07129_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__a21oi_1
X_11553_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04723_ _04728_
+ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10504_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03796_ VGND
+ VGND VPWR VPWR _03811_ sky130_fd_sc_hd__xor2_1
X_14272_ _07070_ _01512_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11484_ _04660_ _04657_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13223_ _05842_ net489 VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10435_ _03747_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13154_ _05998_ _06108_ _06109_ _06110_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__o211a_1
X_10366_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _03675_ VGND
+ VGND VPWR VPWR _03686_ sky130_fd_sc_hd__nand2_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05199_
+ _05129_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__a21o_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _05842_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] VGND
+ VGND VPWR VPWR _06049_ sky130_fd_sc_hd__and2_1
X_10297_ _03625_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _03620_ _03627_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__o211a_1
X_12036_ _05142_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13987_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _06807_ VGND
+ VGND VPWR VPWR _06828_ sky130_fd_sc_hd__nand2_1
X_12938_ _05871_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _05919_ _05920_ _05910_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__o221a_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] VGND VGND VPWR
+ VPWR _05862_ sky130_fd_sc_hd__and3_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ clknet_leaf_46_i_clk _00153_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14539_ clknet_leaf_38_i_clk _00085_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08060_ _01562_ _01656_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08962_ _02321_ net486 _02381_ _02450_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__o211a_1
X_07913_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\] _01521_ _01523_
+ _01453_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__a31o_1
X_08893_ _02389_ _02384_ _02388_ _02369_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07844_ _01465_ net401 VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07775_ net380 net13 _01411_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__mux2_1
X_09514_ _02923_ _02934_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09445_ _02876_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09376_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02813_
+ _02409_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08327_ _01876_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ _01888_ _01890_ _01661_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08258_ _01691_ _01830_ _01689_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08189_ net39 _01329_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__and2_1
X_10220_ _01455_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__clkbuf_4
X_10151_ _03024_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__and2_1
X_10082_ _03442_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__xnor2_1
X_13910_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06716_ VGND
+ VGND VPWR VPWR _06760_ sky130_fd_sc_hd__nand2_1
X_14890_ clknet_leaf_109_i_clk _00435_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13841_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _06700_ _06562_
+ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13772_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06639_
+ _06584_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__o21ai_1
X_10984_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04228_ VGND
+ VGND VPWR VPWR _04229_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12723_ _05733_ _05736_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__and2_1
X_12654_ _05666_ _05672_ _05676_ _05486_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a31o_1
X_15442_ clknet_leaf_27_i_clk _00987_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11605_ _04756_ net161 _04762_ _04768_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12585_ _05609_ _05611_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__nand2_1
X_15373_ clknet_leaf_20_i_clk _00918_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11536_ _04708_ _04705_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__a21o_1
X_14324_ _07113_ _07114_ _06911_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14255_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _07041_ VGND
+ VGND VPWR VPWR _07056_ sky130_fd_sc_hd__xor2_1
X_11467_ _04649_ _04650_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__nand2_1
X_13206_ _06149_ _06151_ _06155_ _05860_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10418_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03732_ VGND
+ VGND VPWR VPWR _03733_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14186_ _06905_ _06994_ _06995_ _06996_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__o211a_1
X_11398_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _04565_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__o41a_1
X_13137_ _05878_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nand2_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND VGND VPWR
+ VPWR _03671_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _06032_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__xnor2_1
X_12019_ _01249_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07560_ diff_valid VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07491_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _01081_ _01085_
+ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09230_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _02685_ _02690_
+ _02691_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09161_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _02629_ VGND
+ VGND VPWR VPWR _02630_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08112_ _01539_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[12\] _01699_ _01705_
+ _01661_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o221a_1
X_09092_ _02559_ _02567_ _02565_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08043_ _01612_ _01620_ _01627_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__a31o_2
XFILLER_0_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09994_ _03352_ _03353_ _03361_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__o21bai_2
X_08945_ _02433_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nor2_1
X_08876_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _02365_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07827_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in VGND VGND VPWR VPWR _01453_
+ sky130_fd_sc_hd__inv_2
X_07758_ net8 net9 _01400_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07689_ net4 _01353_ _01338_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09428_ _02854_ _02858_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09359_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ _05234_ _05435_ _05436_ _05343_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11321_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04520_ VGND
+ VGND VPWR VPWR _04521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14040_ _06563_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06873_
+ _06874_ _06631_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11252_ _04448_ _04452_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _03389_ _03551_ _03552_ _03515_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__o211a_1
X_11183_ _04398_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10134_ _03488_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nor2_1
X_14942_ clknet_leaf_109_i_clk net173 VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10065_ _03426_ _03428_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__xor2_1
X_14873_ clknet_leaf_79_i_clk _00418_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13824_ _06681_ _06684_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10967_ _03997_ net642 _01794_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__o21ai_1
X_13755_ _06625_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _05525_ _05711_
+ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__a21o_1
X_10898_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04152_ VGND
+ VGND VPWR VPWR _04153_ sky130_fd_sc_hd__nand2_1
X_13686_ _06566_ _06567_ _06293_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15425_ clknet_leaf_26_i_clk _00970_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12637_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05641_ VGND
+ VGND VPWR VPWR _05663_ sky130_fd_sc_hd__xor2_2
XFILLER_0_66_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12568_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _05600_ VGND
+ VGND VPWR VPWR _05601_ sky130_fd_sc_hd__and2_1
X_15356_ clknet_leaf_20_i_clk _00901_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11519_ _04680_ _04696_ _04698_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__a21bo_1
X_14307_ _06904_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] VGND
+ VGND VPWR VPWR _07100_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12499_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05541_
+ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15287_ clknet_leaf_17_i_clk _00832_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold207 CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold218 net89 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR net346 sky130_fd_sc_hd__clkdlybuf4s25_1
X_14238_ _07023_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14169_ _06928_ net317 _06981_ _06982_ _06922_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__o221a_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _01881_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _01873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] VGND
+ VGND VPWR VPWR _02188_ sky130_fd_sc_hd__or2_1
X_07612_ _01295_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
X_08592_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[16\] _02125_ VGND VGND VPWR
+ VPWR _02126_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07543_ net407 net317 _01234_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07474_ _01016_ net328 _01198_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ _02657_ _02664_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09144_ _02599_ _02603_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09075_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _02539_ VGND
+ VGND VPWR VPWR _02553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08026_ net36 _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09977_ _03346_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__xor2_1
X_08928_ _02314_ _02418_ _02419_ _02260_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__o211a_1
X_08859_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__or2_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _05000_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _04033_ VGND VGND VPWR
+ VPWR _04083_ sky130_fd_sc_hd__o31a_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10752_ _03669_ _04018_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__nand2_1
X_13540_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _06441_ VGND
+ VGND VPWR VPWR _06442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13471_ _06202_ _06381_ _06382_ _06110_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__o211a_1
X_10683_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03944_ VGND
+ VGND VPWR VPWR _03972_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12422_ _05275_ _05430_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__xnor2_1
X_15210_ clknet_leaf_2_i_clk _00755_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15141_ clknet_leaf_125_i_clk _00686_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12353_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05420_
+ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11304_ _04498_ _04499_ _04505_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15072_ clknet_leaf_118_i_clk _00617_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12284_ _05353_ _05351_ _05356_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14023_ _06850_ _06857_ _06858_ _06569_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__a31o_1
X_11235_ _04378_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11166_ _03619_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__clkbuf_4
X_10117_ _03024_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__and2_1
X_11097_ _04319_ _04311_ _04329_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__and3b_1
X_14925_ clknet_leaf_82_i_clk _00470_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_10048_ _03412_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold90 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
X_14856_ clknet_leaf_79_i_clk _00401_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13807_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _06669_ VGND
+ VGND VPWR VPWR _06670_ sky130_fd_sc_hd__xnor2_1
X_14787_ clknet_leaf_67_i_clk _00332_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_11999_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05081_ VGND
+ VGND VPWR VPWR _05116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13738_ _06610_ _06611_ _06587_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13669_ _06554_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15408_ clknet_leaf_32_i_clk _00953_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15339_ clknet_leaf_48_i_clk _00884_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09900_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _03280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] _03216_
+ _02851_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__o21ai_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _03163_ _03164_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__or2_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _02229_ _02230_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__a21bo_1
X_09693_ _03090_ _03100_ _03101_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08644_ _02015_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _02110_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07526_ _01235_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07457_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _01029_ _01088_
+ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07388_ _01121_ _01126_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09127_ _02156_ _02598_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09058_ _02528_ _02533_ _02536_ _02369_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08009_ net35 _01608_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__and2_1
X_11020_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04251_ _04035_
+ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__o21a_1
X_12971_ _05948_ _03118_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__and2b_1
X_14710_ clknet_leaf_50_i_clk _00255_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11922_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _05047_ VGND
+ VGND VPWR VPWR _05048_ sky130_fd_sc_hd__xnor2_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ clknet_leaf_60_i_clk _00186_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_11853_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _04984_ VGND
+ VGND VPWR VPWR _04985_ sky130_fd_sc_hd__xnor2_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04067_ VGND
+ VGND VPWR VPWR _04068_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11784_ _04923_ _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__nand2_1
X_14572_ clknet_leaf_36_i_clk _00118_ VGND VGND VPWR VPWR diff2\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13523_ _06425_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _06427_ sky130_fd_sc_hd__and2b_1
X_10735_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _04010_ sky130_fd_sc_hd__buf_2
X_10666_ _03945_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _03957_ sky130_fd_sc_hd__and2b_1
X_13454_ _06202_ _06367_ _06368_ _06110_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12405_ _05222_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05465_
+ _05466_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13385_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _06304_ VGND
+ VGND VPWR VPWR _06306_ sky130_fd_sc_hd__nand2_1
X_10597_ _03882_ _03885_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15124_ clknet_leaf_116_i_clk _00669_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_4
X_12336_ _05164_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR out_sintheta[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12267_ _05234_ _05341_ _05342_ _05343_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__o211a_1
X_15055_ clknet_leaf_112_i_clk _00600_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11218_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04428_
+ _04429_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__a21o_1
X_14006_ _06837_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__buf_2
X_12198_ _05282_ _05283_ _05234_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__a21o_1
Xoutput80 net80 VGND VGND VPWR VPWR out_costheta[13] sky130_fd_sc_hd__clkbuf_4
Xoutput91 net91 VGND VGND VPWR VPWR out_costheta[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11149_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__clkbuf_4
X_14908_ clknet_leaf_82_i_clk _00453_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14839_ clknet_leaf_79_i_clk _00384_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08360_ _01915_ _01917_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07311_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _01051_ _01052_
+ _01055_ _01057_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__a221o_1
X_08291_ _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07242_ _00992_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_124_i_clk clknet_4_0_0_i_clk VGND VGND VPWR VPWR clknet_leaf_124_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09814_ _03203_ _03204_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__mux2_1
X_09745_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ _03130_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__nor3_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__or2_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08627_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _02156_ sky130_fd_sc_hd__inv_2
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08558_ _02091_ _02094_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07509_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _01026_ _01223_
+ _01224_ _01030_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__o221a_1
X_08489_ _02011_ _02023_ _02030_ _01924_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10520_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03796_ VGND
+ VGND VPWR VPWR _03825_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10451_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _03762_ VGND
+ VGND VPWR VPWR _03763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13170_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _06112_ VGND
+ VGND VPWR VPWR _06125_ sky130_fd_sc_hd__or2_1
X_10382_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__nor4_1
XFILLER_0_32_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12121_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ _05163_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12052_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05155_
+ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__and2_1
Xhold390 CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] VGND VGND
+ VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _03993_ _04245_ _04246_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__or3_1
X_12954_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__and2b_1
X_11905_ _04771_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _05031_
+ _05032_ _04965_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__o221a_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05874_
+ _05845_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__o21ai_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ clknet_leaf_59_i_clk _00169_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_11836_ _04954_ _04969_ _04970_ _04930_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14555_ clknet_leaf_36_i_clk _00101_ VGND VGND VPWR VPWR diff1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11767_ _04901_ _04902_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__o21ai_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _06352_ VGND
+ VGND VPWR VPWR _06413_ sky130_fd_sc_hd__xnor2_1
X_10718_ net223 _03999_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14486_ clknet_leaf_4_i_clk _00032_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11698_ _04839_ _04840_ _04845_ _04757_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13437_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _06352_ _06347_
+ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer2 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND
+ VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd1_1
X_10649_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ _03920_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nor3_1
XFILLER_0_141_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13368_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _06292_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_41_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15107_ clknet_leaf_111_i_clk _00652_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12319_ _05382_ _05379_ _05388_ _05222_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__a31o_1
XFILLER_0_139_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13299_ _06223_ net577 _06231_ _06233_ _06197_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__o221a_1
X_15038_ clknet_leaf_96_i_clk _00583_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07860_ _01453_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_4
X_07791_ net18 _01423_ net19 VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09530_ _02950_ _02946_ _02953_ _02761_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09461_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _02882_ _02769_
+ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__o21a_1
X_08412_ _01961_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR _01962_ sky130_fd_sc_hd__nor2_1
X_09392_ _02828_ _02832_ _02747_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08343_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] _01897_ _01882_
+ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08274_ _01572_ _01846_ _01847_ _01454_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07989_ _01579_ _01581_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__a21o_1
X_09728_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _03125_ _03121_
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND VGND VPWR VPWR
+ _03134_ sky130_fd_sc_hd__a22o_1
X_09659_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _03070_ VGND
+ VGND VPWR VPWR _03071_ sky130_fd_sc_hd__xnor2_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12670_ _05669_ _05683_ _05681_ _05688_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__and4_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _04776_ _04780_ _04755_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a21o_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14340_ _07127_ _07128_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__or2_1
X_11552_ _04714_ _04716_ _04717_ _04712_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10503_ _03802_ _03810_ _02132_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11483_ _04663_ _04665_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__nand2_1
X_14271_ _06903_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _07068_
+ _07069_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__o2bb2a_1
X_13222_ _05855_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06169_
+ _06170_ _05910_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10434_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03746_ VGND
+ VGND VPWR VPWR _03748_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13153_ _04455_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__clkbuf_4
X_10365_ _03683_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12104_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _05199_
+ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nor2_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _05998_ _06047_ _06048_ _05938_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__o211a_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _03626_ net377 VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12035_ _05139_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13986_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _06807_ VGND
+ VGND VPWR VPWR _06827_ sky130_fd_sc_hd__or2_1
X_12937_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05918_
+ _05842_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _05854_ net635 _05859_ _05861_ _05751_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__o221a_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14607_ clknet_leaf_46_i_clk _00152_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_11819_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04915_ VGND
+ VGND VPWR VPWR _04956_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12799_ _05804_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nor2_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14538_ clknet_leaf_38_i_clk _00084_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14469_ clknet_leaf_5_i_clk _00015_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08961_ _02448_ _02449_ _02322_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__o21ai_1
X_07912_ _01521_ _01523_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[12\]
+ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__a21oi_1
X_08892_ _02384_ _02388_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__a21oi_1
X_07843_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_4
X_07774_ _01416_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09513_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _02938_ VGND
+ VGND VPWR VPWR _02939_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09444_ _02866_ _02868_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__nand2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09375_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08326_ _01877_ _01889_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08257_ _01465_ net630 _01828_ _01833_ _01661_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08188_ _01454_ _01772_ _01775_ _01776_ _01766_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__o311a_1
XFILLER_0_104_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10150_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _03504_ _03185_
+ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__mux2_1
X_10081_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _03410_ VGND
+ VGND VPWR VPWR _03443_ sky130_fd_sc_hd__xnor2_1
X_13840_ _06696_ _06699_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13771_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _06639_
+ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__and2_1
X_10983_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ _04034_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__o21a_1
X_12722_ _05733_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__nor2_1
X_15441_ clknet_leaf_32_i_clk _00986_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ _05666_ _05672_ _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__a21oi_1
X_11604_ _04758_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15372_ clknet_leaf_20_i_clk _00917_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12584_ _05501_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14323_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__nor2_1
X_11535_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _04692_ VGND
+ VGND VPWR VPWR _04713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14254_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[4\]
+ _07041_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__o41a_1
XFILLER_0_150_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11466_ _04646_ _04648_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13205_ _06149_ _06151_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10417_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _03650_ _03720_
+ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11397_ _04570_ _04574_ _04581_ _04586_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__and4b_1
X_14185_ _04455_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13136_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__or4_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _03623_ _03668_ _03670_ _03515_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__o211a_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _06025_ _06029_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__o21ai_1
X_10279_ _03607_ net266 _03568_ _03615_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__o211a_1
X_12018_ _05130_ net183 _04979_ _05131_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13969_ _06732_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND
+ VGND VPWR VPWR _06813_ sky130_fd_sc_hd__or2_1
X_07490_ _01016_ net255 _01210_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09160_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _02628_ VGND
+ VGND VPWR VPWR _02629_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08111_ _01556_ _01704_ _01480_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09091_ _02559_ _02565_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08042_ net35 net53 _01627_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__a31o_1
X_09993_ _03184_ _03362_ _03363_ _03292_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08944_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02432_ VGND
+ VGND VPWR VPWR _02434_ sky130_fd_sc_hd__nor2_1
X_08875_ _02329_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _02374_ _02375_ _02309_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__o221a_1
X_07826_ _01452_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
X_07757_ _01404_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07688_ net4 _01353_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09427_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _02857_ VGND
+ VGND VPWR VPWR _02861_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09358_ _02750_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08309_ _01867_ net164 _01823_ _01875_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _02745_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11320_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04519_ VGND
+ VGND VPWR VPWR _04520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11251_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _04451_ VGND
+ VGND VPWR VPWR _04457_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10202_ _03190_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND
+ VGND VPWR VPWR _03552_ sky130_fd_sc_hd__or2_1
X_11182_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND VPWR
+ VPWR _04399_ sky130_fd_sc_hd__a21oi_1
X_10133_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03486_ VGND
+ VGND VPWR VPWR _03489_ sky130_fd_sc_hd__nor2_1
X_14941_ clknet_leaf_109_i_clk net180 VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10064_ _03427_ _03422_ _03418_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14872_ clknet_leaf_79_i_clk _00417_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_13823_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] _06681_ _06684_
+ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13754_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _06615_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__and3_1
X_10966_ _04203_ _04209_ _04212_ _03997_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12705_ _05721_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
X_13685_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__or2_1
X_10897_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04151_ VGND
+ VGND VPWR VPWR _04152_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15424_ clknet_leaf_25_i_clk _00969_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12636_ _05662_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15355_ clknet_leaf_19_i_clk _00900_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12567_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05599_ VGND
+ VGND VPWR VPWR _05600_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14306_ _07059_ _07098_ _07099_ _06996_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__o211a_1
X_11518_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04684_ _04697_
+ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__o21ai_1
X_15286_ clknet_leaf_51_i_clk _00831_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12498_ _05203_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _05535_ _05540_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__o31a_1
Xhold208 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR
+ VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND VGND
+ VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ _07029_ _07039_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__and2b_1
X_11449_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _04634_ VGND
+ VGND VPWR VPWR _04635_ sky130_fd_sc_hd__xor2_2
XFILLER_0_150_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14168_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06980_
+ _01862_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__o21ai_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _06069_ _06078_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__and2_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _06647_ _06917_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__nand2_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08660_ _02185_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07611_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\] _01294_ _01282_ VGND
+ VGND VPWR VPWR _01295_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_6_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_6_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_08591_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[17\] _02122_ _02124_ VGND
+ VGND VPWR VPWR _02125_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07542_ _01243_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
X_07473_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _01159_ _01196_
+ _01197_ _01030_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__o221a_1
X_09212_ _02655_ _02662_ _02663_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09143_ _02613_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09074_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02541_ VGND
+ VGND VPWR VPWR _02552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08025_ net54 VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09976_ _03334_ _03338_ _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08927_ _02315_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _02419_ sky130_fd_sc_hd__or2_1
X_08858_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _02360_
+ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__xor2_1
X_07809_ _01440_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[16\] _02299_ VGND VGND VPWR
+ VPWR _02304_ sky130_fd_sc_hd__and2_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _04082_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10751_ _04010_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13470_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND
+ VGND VPWR VPWR _06382_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10682_ _03971_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12421_ _05480_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15140_ clknet_leaf_125_i_clk _00685_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_12352_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _05404_ VGND
+ VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11303_ _04503_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15071_ clknet_leaf_102_i_clk _00616_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12283_ _05353_ _05351_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14022_ _06850_ _06857_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__a21oi_1
X_11234_ net422 _04438_ _04437_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a21oi_1
X_11165_ _04377_ net260 _04219_ _04386_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10116_ _03472_ _03473_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ _03182_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a2bb2o_1
X_11096_ _04012_ net621 _04330_ _04331_ _04059_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14924_ clknet_leaf_82_i_clk _00469_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10047_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _03410_ _03411_
+ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__and3_1
Xhold80 net97 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net111 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14855_ clknet_leaf_79_i_clk _00400_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13806_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _06586_ VGND VGND
+ VPWR VPWR _06669_ sky130_fd_sc_hd__o31a_1
XFILLER_0_98_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14786_ clknet_leaf_67_i_clk _00331_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11998_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _05081_ VGND
+ VGND VPWR VPWR _05115_ sky130_fd_sc_hd__or2_1
X_13737_ _06610_ _06605_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__nand2_1
X_10949_ _04189_ _04194_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13668_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15407_ clknet_leaf_32_i_clk _00952_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12619_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _05641_ VGND
+ VGND VPWR VPWR _05647_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13599_ _06486_ _06487_ _06491_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15338_ clknet_leaf_49_i_clk _00883_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_130_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15269_ clknet_leaf_12_i_clk _00814_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09830_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _03204_ VGND VGND
+ VPWR VPWR _03221_ sky130_fd_sc_hd__and4_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03151_ VGND
+ VGND VPWR VPWR _03164_ sky130_fd_sc_hd__nor2_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[10\] _02233_ VGND VGND VPWR
+ VPWR _02234_ sky130_fd_sc_hd__xnor2_1
X_09692_ _02891_ _03089_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__or2_1
X_08643_ _01879_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _01981_ _02109_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__and2_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ net373 net316 _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07456_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _01081_ _01184_
+ _01085_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07387_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _01017_ _01122_
+ _01125_ _01072_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09126_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] _02597_ VGND
+ VGND VPWR VPWR _02598_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ _02528_ _02533_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ net53 VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09959_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _03331_ VGND
+ VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xnor2_1
X_12970_ _05860_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _05946_
+ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__a22oi_1
X_11921_ _05046_ _04952_ net114 CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__a31o_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ clknet_leaf_60_i_clk _00185_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11852_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _04983_ VGND
+ VGND VPWR VPWR _04984_ sky130_fd_sc_hd__xnor2_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ clknet_leaf_36_i_clk _00117_ VGND VGND VPWR VPWR diff2\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04915_ VGND
+ VGND VPWR VPWR _04924_ sky130_fd_sc_hd__or2_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13522_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _06425_ VGND
+ VGND VPWR VPWR _06426_ sky130_fd_sc_hd__and2b_1
X_10734_ _03995_ net158 _04003_ _04009_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13453_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _06368_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10665_ _03954_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12404_ _05464_ _05460_ _05461_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__o31a_1
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13384_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _06304_ VGND
+ VGND VPWR VPWR _06305_ sky130_fd_sc_hd__nor2_1
X_10596_ _03891_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__or2_1
X_15123_ clknet_leaf_116_i_clk _00668_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12335_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05375_ VGND VGND
+ VPWR VPWR _05404_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15054_ clknet_leaf_112_i_clk net139 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12266_ _04455_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14005_ _06842_ _06843_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11217_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] _04428_
+ _04378_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__o21ai_1
X_12197_ _05281_ _05272_ _05274_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__nand3_1
Xoutput70 net70 VGND VGND VPWR VPWR out_alpha[4] sky130_fd_sc_hd__clkbuf_4
Xoutput81 net81 VGND VGND VPWR VPWR out_costheta[14] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 VGND VGND VPWR VPWR out_costheta[8] sky130_fd_sc_hd__clkbuf_4
X_11148_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11079_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__inv_2
X_14907_ clknet_leaf_82_i_clk _00452_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14838_ clknet_leaf_75_i_clk _00383_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14769_ clknet_leaf_52_i_clk _00314_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07310_ _01056_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08290_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _01861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07241_ _00999_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09813_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__clkbuf_4
X_09744_ _02754_ net429 _03017_ _03148_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__o211a_1
X_09675_ _02755_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03084_
+ _03085_ _03013_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__o221a_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _02155_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _02092_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07508_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _01122_ _01167_
+ _01046_ _01072_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__a221o_1
X_08488_ _02011_ _02023_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07439_ _01171_ _01165_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10450_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03761_ VGND
+ VGND VPWR VPWR _03762_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09109_ _02576_ _02581_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10381_ _03694_ _03695_ _03692_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__a21o_1
X_12120_ _05130_ _05211_ _05212_ _05080_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12051_ _04829_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _05145_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__o31a_1
Xhold380 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold391 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR VPWR
+ net508 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ _04238_ _04231_ _04244_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12953_ _05871_ net492 _05931_ _05932_ _05910_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11904_ _05018_ _05021_ _05030_ _04758_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12884_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _05874_
+ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and2_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ clknet_leaf_60_i_clk _00168_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11835_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__or4_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ clknet_leaf_34_i_clk _00100_ VGND VGND VPWR VPWR diff1\[13\] sky130_fd_sc_hd__dfxtp_1
X_11766_ _04907_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _06352_ _06410_ _06411_ _06385_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__o2bb2a_1
X_10717_ _03995_ net240 _03620_ _04000_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14485_ clknet_leaf_24_i_clk _00031_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_1
X_11697_ _04839_ _04840_ _04845_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13436_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__clkbuf_4
X_10648_ _03606_ _03939_ _03940_ _03780_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__o211a_1
Xrebuffer3 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] VGND VGND
+ VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _06287_
+ _06286_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__a21oi_1
X_10579_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03871_ VGND
+ VGND VPWR VPWR _03877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15106_ clknet_leaf_111_i_clk net219 VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12318_ _05382_ _05379_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13298_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _06230_
+ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15037_ clknet_leaf_101_i_clk _00582_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12249_ _05326_ _05327_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07790_ _01426_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09460_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] VGND VGND VPWR
+ VPWR _02891_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08411_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[1\] VGND VGND VPWR VPWR
+ _01961_ sky130_fd_sc_hd__inv_2
X_09391_ _02829_ _02831_ _02772_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__mux2_1
X_08342_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] _01898_ _01882_
+ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08273_ _01572_ _01743_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07988_ net32 net50 VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__and2_1
X_09727_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03132_ VGND
+ VGND VPWR VPWR _03133_ sky130_fd_sc_hd__xor2_2
X_09658_ _02770_ _03069_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__and2_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\] _02139_ VGND VGND VPWR
+ VPWR _02140_ sky130_fd_sc_hd__xnor2_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _03008_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _04776_ _04780_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__nor2_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11551_ _04396_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND
+ VGND VPWR VPWR _04727_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ _03642_ _03808_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__and3_1
X_14270_ _07067_ _07065_ _07066_ _06902_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__a31o_1
X_11482_ _04664_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13221_ _06159_ _06165_ _06168_ _05860_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__a31o_1
X_10433_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _03746_ VGND
+ VGND VPWR VPWR _03747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13152_ _05853_ net539 VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10364_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _03682_ VGND
+ VGND VPWR VPWR _03684_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ _05197_ _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__or2b_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND
+ VGND VPWR VPWR _06048_ sky130_fd_sc_hd__or2_1
X_10295_ _03608_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__clkbuf_4
X_12034_ _03619_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__buf_4
X_13985_ _06826_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
X_12936_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05918_
+ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12867_ _05567_ _05857_ _05858_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__a31o_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_123_i_clk clknet_4_0_0_i_clk VGND VGND VPWR VPWR clknet_leaf_123_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11818_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _04930_ VGND
+ VGND VPWR VPWR _04955_ sky130_fd_sc_hd__nor2_1
X_14606_ clknet_leaf_47_i_clk _00151_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12798_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05781_ VGND
+ VGND VPWR VPWR _05805_ sky130_fd_sc_hd__and2_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ clknet_leaf_38_i_clk _00083_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_11749_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04794_ _04884_
+ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14468_ clknet_leaf_4_i_clk _00014_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13419_ _06336_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__buf_2
X_14399_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _07157_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08960_ _02433_ _02440_ _02447_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__nor3_1
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07911_ _01328_ _01522_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__nand2_1
X_08891_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR _02389_ sky130_fd_sc_hd__inv_2
X_07842_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.valid_in VGND VGND VPWR VPWR _01464_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07773_ net360 net12 _01411_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__mux2_1
X_09512_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _02937_ VGND
+ VGND VPWR VPWR _02938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09443_ _02874_ _02875_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__nor2_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09374_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ _02806_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _02817_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_19_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08325_ _01886_ _01887_ _01550_ _01883_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08256_ _01831_ _01832_ _01529_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08187_ _01464_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[17\] VGND VGND VPWR
+ VPWR _01776_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10080_ _03431_ _03438_ _03432_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13770_ _06293_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _06632_ _06638_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__o31a_1
X_10982_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND VGND VPWR
+ VPWR _04227_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_40_i_clk clknet_4_11_0_i_clk VGND VGND VPWR VPWR clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12721_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _05735_ VGND
+ VGND VPWR VPWR _05736_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15440_ clknet_leaf_27_i_clk _00985_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12652_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _05641_ VGND
+ VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xor2_1
X_11603_ _04756_ net138 _04762_ _04767_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__o211a_1
X_15371_ clknet_leaf_20_i_clk _00916_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12583_ net586 VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_55_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14322_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__and2_1
X_11534_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _04692_ VGND
+ VGND VPWR VPWR _04712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14253_ _07029_ _07046_ _07039_ _07051_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__and4b_1
X_11465_ _04646_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13204_ _05930_ _06136_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10416_ _03731_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14184_ _06907_ net432 VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__or2_1
X_11396_ _04431_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04587_
+ _04588_ _04539_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__o221a_1
XFILLER_0_110_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13135_ _06085_ _06089_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10347_ _03621_ _03669_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _06010_ VGND
+ VGND VPWR VPWR _06033_ sky130_fd_sc_hd__nand2_1
X_10278_ net265 _03609_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__or2_1
X_12017_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] _01250_
+ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13968_ _06804_ _06811_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12919_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _05890_ VGND
+ VGND VPWR VPWR _05904_ sky130_fd_sc_hd__or4_1
X_13899_ _06748_ _06749_ _06750_ _06553_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08110_ _01691_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09090_ _02542_ _02547_ _02566_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08041_ net36 net54 VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_i_clk clknet_0_i_clk VGND VGND VPWR VPWR clknet_4_2_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09992_ _03290_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _03363_ sky130_fd_sc_hd__or2_1
X_08943_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02432_ VGND
+ VGND VPWR VPWR _02433_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08874_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02373_
+ _02320_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__o21ai_1
X_07825_ net502 _01451_ _00992_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07756_ net472 _01403_ _01358_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__mux2_1
X_07687_ _01353_ _01354_ net227 _01333_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_149_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09426_ _02748_ _02859_ _02860_ _02260_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09357_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _02802_
+ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08308_ _01870_ net650 VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _02744_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08239_ _01636_ _01670_ _01652_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11250_ _04442_ _04453_ _04454_ _04456_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10201_ _03548_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11181_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND VPWR
+ VPWR _04398_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10132_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14940_ clknet_leaf_110_i_clk net235 VGND VGND VPWR VPWR CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10063_ _03420_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__inv_2
X_14871_ clknet_leaf_78_i_clk _00416_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_13822_ _06683_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13753_ _06561_ net561 _06485_ _06624_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__o211a_1
X_10965_ _04203_ _04209_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__o21ai_1
X_12704_ _05652_ _05720_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__and2_1
X_13684_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10896_ _04034_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__and2_1
X_12635_ _05652_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__and2_1
X_15423_ clknet_leaf_26_i_clk _00968_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15354_ clknet_leaf_29_i_clk _00899_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12566_ _05526_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11517_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _04684_ _04674_
+ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14305_ _06909_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND
+ VGND VPWR VPWR _07099_ sky130_fd_sc_hd__or2_1
X_15285_ clknet_leaf_16_i_clk _00830_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12497_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05539_
+ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14236_ _07032_ _07035_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__nor2_1
Xhold209 diff1\[8\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _04633_ VGND
+ VGND VPWR VPWR _04634_ sky130_fd_sc_hd__xor2_2
XFILLER_0_33_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14167_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06980_
+ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04545_ VGND
+ VGND VPWR VPWR _04574_ sky130_fd_sc_hd__xnor2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _05844_ _06075_ _06076_ _06077_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__a31o_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _06910_ net323 _06920_ _06921_ _06922_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__o221a_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _06017_ _06015_ _06016_ _05860_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07610_ r_i_alpha1\[8\] _01293_ _01276_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__mux2_1
X_08590_ _02123_ _01549_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[17\] VGND
+ VGND VPWR VPWR _02124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07541_ net366 net320 _01234_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07472_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _01122_ _01092_
+ _01047_ _01072_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__a221o_1
X_09211_ _02674_ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09142_ _02611_ _02612_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09073_ _02551_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08024_ _01463_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\] _01460_ _01623_
+ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09975_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03332_ VGND
+ VGND VPWR VPWR _03347_ sky130_fd_sc_hd__nand2_1
X_08926_ _02412_ _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08857_ _01959_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ _02355_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__o22a_1
X_07808_ net383 _01439_ _01411_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _02290_ _02303_ _02132_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__o21a_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07739_ _01338_ _01391_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__nand2_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10750_ _04011_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _04021_ _04022_ _03814_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09409_ net440 VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10681_ _03535_ _03970_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ _05290_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12351_ _05366_ _05370_ _05410_ _05417_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11302_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04502_ VGND
+ VGND VPWR VPWR _04504_ sky130_fd_sc_hd__or2_1
X_15070_ clknet_leaf_102_i_clk _00615_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12282_ _04996_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14021_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _06837_ VGND
+ VGND VPWR VPWR _06858_ sky130_fd_sc_hd__xor2_1
X_11233_ _04376_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11164_ net138 _04379_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__or2_1
X_10115_ _03469_ _03471_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__nor2_1
X_11095_ _04317_ _04320_ _04329_ _04047_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a31o_1
X_14923_ clknet_leaf_82_i_clk _00468_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_10046_ _03410_ _03411_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold70 _00483_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 diff3\[10\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ clknet_leaf_79_i_clk _00399_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13805_ _06668_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
X_11997_ _04771_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05113_
+ _05114_ _04965_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__o221a_1
X_14785_ clknet_leaf_70_i_clk _00330_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10948_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04177_ VGND
+ VGND VPWR VPWR _04198_ sky130_fd_sc_hd__xnor2_1
X_13736_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND
+ VPWR VPWR _06610_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10879_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04134_ VGND
+ VGND VPWR VPWR _04136_ sky130_fd_sc_hd__or2_1
X_13667_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _06553_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15406_ clknet_leaf_32_i_clk _00951_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12618_ _05632_ _05645_ _05646_ _05343_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13598_ _06210_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _06485_
+ _06494_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12549_ _05581_ _05583_ _05485_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15337_ clknet_leaf_49_i_clk _00882_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15268_ clknet_leaf_10_i_clk _00813_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14219_ _07022_ _07024_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15199_ clknet_leaf_1_i_clk _00744_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09760_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _03151_ VGND
+ VGND VPWR VPWR _03163_ sky130_fd_sc_hd__and2_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[11\] _02232_ VGND VGND VPWR
+ VPWR _02233_ sky130_fd_sc_hd__xor2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _03054_ _03063_ _03074_ _03083_ _03093_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_83_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08642_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[4\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[3\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[2\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\]
+ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__or4_4
XFILLER_0_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08573_ _01865_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02107_
+ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__a22o_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07524_ _01012_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07455_ _01051_ _01048_ _01049_ _01076_ _01055_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07386_ _01123_ _01124_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__and2_1
X_09125_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _02341_ VGND VGND VPWR
+ VPWR _02597_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09056_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _02535_ VGND
+ VGND VPWR VPWR _02536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08007_ _01463_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[5\] _01460_ _01607_
+ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09958_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ _03315_ _03205_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__o31a_1
X_08909_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _02399_
+ _02344_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__o21ai_1
X_09889_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] VGND VGND
+ VPWR VPWR _03271_ sky130_fd_sc_hd__inv_2
X_11920_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] VGND VGND VPWR
+ VPWR _05046_ sky130_fd_sc_hd__inv_2
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__and2b_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _04023_ net400 _04065_ _04066_ _04059_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__o221a_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ clknet_leaf_34_i_clk _00116_ VGND VGND VPWR VPWR diff2\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _04915_ VGND
+ VGND VPWR VPWR _04923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10733_ _03997_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\]
+ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__or2_1
X_13521_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06424_ VGND
+ VGND VPWR VPWR _06425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13452_ _06365_ _06366_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__nor2_1
X_10664_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03944_ VGND
+ VGND VPWR VPWR _03955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12403_ _05460_ _05461_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_91_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13383_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _06303_ VGND
+ VGND VPWR VPWR _06304_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10595_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03890_ VGND
+ VGND VPWR VPWR _03892_ sky130_fd_sc_hd__nor2_1
X_15122_ clknet_leaf_116_i_clk _00667_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR
+ VPWR _05403_ sky130_fd_sc_hd__inv_2
X_15053_ clknet_leaf_112_i_clk net135 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12265_ _05139_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _05342_ sky130_fd_sc_hd__or2_1
X_14004_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06837_ VGND
+ VGND VPWR VPWR _06843_ sky130_fd_sc_hd__nand2_1
X_11216_ _04426_ _04427_ _04414_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__mux2_1
X_12196_ _05272_ _05274_ _05281_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__a21o_1
Xoutput60 net60 VGND VGND VPWR VPWR out_alpha[11] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 VGND VGND VPWR VPWR out_alpha[5] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 VGND VGND VPWR VPWR out_costheta[15] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 VGND VGND VPWR VPWR out_costheta[9] sky130_fd_sc_hd__clkbuf_4
X_11147_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11078_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04314_ VGND
+ VGND VPWR VPWR _04315_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14906_ clknet_leaf_82_i_clk _00451_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10029_ _03394_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14837_ clknet_leaf_77_i_clk _00382_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14768_ clknet_leaf_52_i_clk _00313_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13719_ _06593_ _06595_ _06587_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14699_ clknet_leaf_63_i_clk _00244_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07240_ net329 net20 _00993_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09812_ _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__buf_2
X_09743_ _03143_ _03146_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09674_ _03072_ _03075_ _03083_ _02746_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__a31o_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _01981_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__and2_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[13\] _02083_ _01881_ VGND
+ VGND VPWR VPWR _02093_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07507_ _01022_ _01163_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08487_ _02028_ _02029_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__and2_2
XFILLER_0_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07438_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] VGND VGND
+ VPWR VPWR _01171_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07369_ _01108_ _01109_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09108_ _02576_ _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10380_ _03698_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09039_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] VGND VGND VPWR
+ VPWR _02520_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12050_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] _05148_
+ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__nand2_1
Xhold370 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] VGND VGND
+ VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR
+ VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND
+ VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _04238_ _04231_ _04244_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__and3_1
X_12952_ _05930_ net471 _05842_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__a21o_1
X_11903_ _05018_ _05021_ _05030_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__o21a_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _05872_ _05873_ _05566_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__mux2_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ clknet_leaf_60_i_clk _00167_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_11834_ _04957_ _04962_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__or2_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11765_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04906_ VGND
+ VGND VPWR VPWR _04908_ sky130_fd_sc_hd__or2_1
X_14553_ clknet_leaf_34_i_clk _00099_ VGND VGND VPWR VPWR diff1\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10716_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] _03999_
+ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__or2_1
X_13504_ _06396_ _06399_ _06406_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11696_ _04843_ _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14484_ clknet_leaf_25_i_clk _00030_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10647_ _03608_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND
+ VGND VPWR VPWR _03940_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13435_ _06337_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer4 _05236_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_1
X_13366_ _06223_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ _06289_ _06290_ _06285_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__o221a_1
X_10578_ _03626_ net405 _03875_ _03876_ _03814_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__o221a_1
X_15105_ clknet_leaf_111_i_clk net184 VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12317_ _05386_ _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13297_ _06204_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12248_ _05319_ _05322_ _05318_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__o21ai_1
X_15036_ clknet_leaf_92_i_clk _00581_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12179_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _05254_ _05256_
+ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08410_ _01867_ _01957_ _01960_ _01552_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__o211a_1
X_09390_ _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08341_ _01876_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ _01823_ _01902_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08272_ _01738_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07987_ _01587_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__nand2_4
X_09726_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03131_ VGND
+ VGND VPWR VPWR _03132_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09657_ _03048_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__or2_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[1\]
+ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__and2b_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _02497_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__and2_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08539_ _02065_ _02073_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11550_ _04376_ _04725_ _04726_ _04456_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10501_ _03807_ _03803_ _03804_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_80_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11481_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04662_ VGND
+ VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nor2_1
X_13220_ _06159_ _06165_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10432_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03745_ VGND
+ VGND VPWR VPWR _03746_ sky130_fd_sc_hd__xor2_1
X_13151_ _06105_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10363_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _03682_ VGND
+ VGND VPWR VPWR _03683_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12102_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05192_
+ _05164_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a21o_1
X_13082_ _06044_ _06046_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__xnor2_1
X_10294_ _03608_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__buf_2
X_12033_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13984_ _01253_ _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__and2_1
X_12935_ _05916_ _05917_ _05878_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _05841_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__clkbuf_4
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ clknet_leaf_47_i_clk _00150_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11817_ _04941_ _04944_ _04948_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__or3_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _05781_ VGND
+ VGND VPWR VPWR _05804_ sky130_fd_sc_hd__nor2_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ clknet_leaf_38_i_clk _00082_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11748_ _04892_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14467_ clknet_leaf_39_i_clk _00013_ VGND VGND VPWR VPWR r_i_alpha1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11679_ _04756_ _04828_ _04830_ _04739_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13418_ _06332_ _06334_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14398_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _07157_ _07172_
+ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__o21a_1
X_13349_ _06274_ _06275_ _06235_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15019_ clknet_leaf_98_i_clk _00564_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_07910_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[11\] _01515_ VGND VGND
+ VPWR VPWR _01522_ sky130_fd_sc_hd__or2_1
X_08890_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _02382_
+ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__or2_1
X_07841_ _01457_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07772_ _01415_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
X_09511_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ _02918_ _02771_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__o31a_1
XFILLER_0_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09442_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02873_ VGND
+ VGND VPWR VPWR _02875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09373_ _02757_ net530 _02815_ _02816_ _02689_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08324_ _01550_ _01883_ _01886_ _01887_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08255_ _01691_ _01830_ _01470_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08186_ _01773_ _01774_ _01330_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09709_ _03105_ _03116_ _02750_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__mux2_1
X_10981_ _04221_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] VGND
+ VGND VPWR VPWR _04226_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12720_ _05525_ _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12651_ _05632_ _05673_ _05674_ _05675_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11602_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _04765_
+ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or2_1
X_12582_ _05521_ net352 _05612_ _05613_ _05544_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__o221a_1
X_15370_ clknet_leaf_21_i_clk _00915_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14321_ _07059_ _07111_ _07112_ _01475_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11533_ _04391_ net520 _04710_ _04711_ _04539_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11464_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _04647_ VGND
+ VGND VPWR VPWR _04648_ sky130_fd_sc_hd__xnor2_1
X_14252_ _06911_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _07052_
+ _07053_ _01456_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13203_ _06154_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_1
X_10415_ _03535_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11395_ _04579_ _04582_ _04586_ _04396_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__a31o_1
X_14183_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _06993_
+ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10346_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _03669_ sky130_fd_sc_hd__buf_2
X_13134_ _06092_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] _06003_ VGND
+ VGND VPWR VPWR _06032_ sky130_fd_sc_hd__xnor2_1
X_10277_ _03607_ net130 _03568_ _03614_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__o211a_1
X_12016_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13967_ _06809_ _06810_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_88_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12918_ _05871_ net557 _05902_ _05903_ _05751_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13898_ _06736_ _06740_ _06743_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _05844_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__buf_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14519_ clknet_leaf_32_i_clk _00065_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08040_ _01636_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__nand2_4
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09991_ _03354_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08942_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _02431_ VGND
+ VGND VPWR VPWR _02432_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08873_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02373_
+ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07824_ net11 _01449_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07755_ net8 _01400_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07686_ net20 _01350_ _01345_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09425_ _02804_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _02860_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ _02800_ _02801_ _02772_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08307_ _01867_ net165 _01823_ _01874_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09287_ _02320_ _02310_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08238_ _01717_ net458 _01635_ _01817_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08169_ _01750_ _01738_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10200_ _03539_ _03542_ _03549_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11180_ _04390_ net506 _04395_ _04397_ _04360_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__o221a_1
X_10131_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _03486_ VGND
+ VGND VPWR VPWR _03487_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_122_i_clk clknet_4_0_0_i_clk VGND VGND VPWR VPWR clknet_leaf_122_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10062_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03410_ VGND
+ VGND VPWR VPWR _03426_ sky130_fd_sc_hd__xor2_1
X_14870_ clknet_leaf_84_i_clk _00415_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_13821_ _06682_ _06586_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13752_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06622_
+ _06623_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__a21o_1
X_10964_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _04177_ VGND
+ VGND VPWR VPWR _04212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12703_ _05486_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _05718_
+ _05719_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13683_ _06562_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__clkbuf_4
X_10895_ _04108_ _04149_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15422_ clknet_leaf_25_i_clk _00967_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12634_ _05489_ _05658_ _05659_ _05660_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15353_ clknet_leaf_48_i_clk _00898_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12565_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__or4_2
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14304_ _07096_ _07097_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__xnor2_1
X_11516_ _04676_ _04685_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15284_ clknet_leaf_16_i_clk _00829_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12496_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\]
+ _05528_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14235_ _06905_ _07037_ _07038_ _06996_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11447_ _04412_ net652 VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11378_ _04442_ _04572_ _04573_ _04456_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__o211a_1
X_14166_ _06647_ _06977_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__o21a_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _05841_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] VGND
+ VGND VPWR VPWR _06077_ sky130_fd_sc_hd__and2_1
X_10329_ _03652_ _03653_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__a21oi_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _01474_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__clkbuf_4
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _06015_ _06016_ _06017_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14999_ clknet_leaf_108_i_clk _00544_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_07540_ _01242_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07471_ _01022_ _01090_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09210_ _02237_ _02673_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09141_ _02607_ _02610_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09072_ _02497_ _02550_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08023_ _01330_ _01617_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09974_ _03344_ _03345_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08925_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _02416_ VGND
+ VGND VPWR VPWR _02417_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_54_i_clk clknet_4_14_0_i_clk VGND VGND VPWR VPWR clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08856_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _02348_
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] VGND VGND VPWR
+ VPWR _02359_ sky130_fd_sc_hd__a21oi_1
X_07807_ _01003_ _01435_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__xnor2_1
X_08787_ _02301_ _02302_ _01873_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__and3b_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ net19 _01385_ net20 VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__a21o_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07669_ net228 _01333_ _01337_ _01340_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09408_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _02829_ _02772_
+ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__a41o_1
X_10680_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _03969_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09339_ _02757_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _02786_ _02787_ _02689_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__o221a_1
XFILLER_0_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12350_ _05407_ _05408_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11301_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04502_ VGND
+ VGND VPWR VPWR _04503_ sky130_fd_sc_hd__nand2_1
X_12281_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _05354_ VGND
+ VGND VPWR VPWR _05355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11232_ _04377_ _04440_ _04441_ _04063_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14020_ _06853_ _06851_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__or2b_1
X_11163_ _04377_ net261 _04219_ _04385_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10114_ _03469_ _03471_ _03182_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__a21o_1
X_11094_ _04317_ _04320_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a21oi_1
X_14922_ clknet_leaf_88_i_clk _00467_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_10045_ _03407_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03391_
+ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 net100 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold71 diff1\[14\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 diff2\[8\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ clknet_leaf_79_i_clk _00398_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold93 CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND VGND
+ VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _06667_ _01512_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__and2b_1
X_14784_ clknet_leaf_70_i_clk _00329_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11996_ _05111_ _05112_ _04786_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13735_ _06565_ net576 _06608_ _06609_ _06526_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__o221a_1
X_10947_ _04048_ _04196_ _04197_ _04063_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13666_ _06552_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
X_10878_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04134_ VGND
+ VGND VPWR VPWR _04135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15405_ clknet_leaf_32_i_clk _00950_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12617_ _05492_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] VGND
+ VGND VPWR VPWR _05646_ sky130_fd_sc_hd__or2_1
X_13597_ _06492_ _06493_ _06232_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15336_ clknet_leaf_38_i_clk _00881_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12548_ _05570_ _05574_ _05582_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15267_ clknet_leaf_10_i_clk _00812_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12479_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _05525_ sky130_fd_sc_hd__inv_2
X_14218_ _07019_ _07023_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[3\]
+ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__a21oi_1
X_15198_ clknet_leaf_0_i_clk _00743_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14149_ _06928_ net322 _06964_ _06965_ _06922_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _01881_ _02231_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__nand2_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _03098_ VGND
+ VGND VPWR VPWR _03099_ sky130_fd_sc_hd__xnor2_1
X_08641_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR VPWR
+ _02169_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08572_ _02103_ _02106_ _01868_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__o21a_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07523_ net304 VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07454_ _01095_ net617 _01182_ _01183_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07385_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _01108_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09124_ _02152_ _02587_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09055_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _02534_ VGND
+ VGND VPWR VPWR _02535_ sky130_fd_sc_hd__xor2_2
XFILLER_0_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08006_ _01465_ _01606_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__nand2_1
Xhold530 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09957_ _03189_ net441 _03017_ _03330_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__o211a_1
X_08908_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _02402_ _02403_ _02309_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o221a_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _03237_ net541 _03269_ _03270_ _03258_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08839_ _02344_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__or2_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _04769_ net271 _04979_ _04982_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__o211a_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _04064_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] _03994_
+ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__a21o_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _04769_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _04762_
+ _04922_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__o211a_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13520_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__and2b_1
X_10732_ _03995_ net172 _04003_ _04008_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13451_ _06364_ _06356_ _06361_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10663_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _03944_ VGND
+ VGND VPWR VPWR _03954_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12402_ _05462_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10594_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03890_ VGND
+ VGND VPWR VPWR _03891_ sky130_fd_sc_hd__and2_1
X_13382_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[12\]
+ _06235_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15121_ clknet_leaf_116_i_clk _00666_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12333_ _05402_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15052_ clknet_leaf_111_i_clk _00597_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12264_ _05339_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14003_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _06807_ VGND
+ VGND VPWR VPWR _06842_ sky130_fd_sc_hd__or2_1
X_11215_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _04421_
+ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__or2_1
X_12195_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _05280_ VGND
+ VGND VPWR VPWR _05281_ sky130_fd_sc_hd__xnor2_1
Xoutput61 net61 VGND VGND VPWR VPWR out_alpha[12] sky130_fd_sc_hd__clkbuf_4
Xoutput72 net72 VGND VGND VPWR VPWR out_alpha[6] sky130_fd_sc_hd__clkbuf_4
X_11146_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _04374_ sky130_fd_sc_hd__inv_2
Xoutput83 net83 VGND VGND VPWR VPWR out_costheta[16] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 VGND VGND VPWR VPWR out_sintheta[0] sky130_fd_sc_hd__clkbuf_4
X_11077_ _04035_ _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__nand2_1
X_14905_ clknet_leaf_82_i_clk _00450_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10028_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03393_ VGND
+ VGND VPWR VPWR _03395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14836_ clknet_leaf_77_i_clk _00381_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14767_ clknet_leaf_52_i_clk _00312_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11979_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _05072_ VGND
+ VGND VPWR VPWR _05099_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13718_ _06594_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14698_ clknet_leaf_61_i_clk _00243_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13649_ _06211_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _06537_
+ _06538_ _06526_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15319_ clknet_leaf_22_i_clk _00864_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09811_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _03205_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09742_ _03143_ _03146_ _02750_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09673_ _03072_ _03075_ _03083_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a21oi_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _01869_ _02150_ _02151_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[14\] VGND VGND VPWR VPWR
+ _02092_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07506_ _01016_ net214 _01222_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08486_ _02024_ _02027_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07437_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _01161_ VGND
+ VGND VPWR VPWR _01170_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _01099_ VGND
+ VGND VPWR VPWR _01109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09107_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[1\] _02580_ VGND
+ VGND VPWR VPWR _02581_ sky130_fd_sc_hd__xnor2_1
X_07299_ _01017_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\]
+ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09038_ _02507_ _02516_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold360 net81 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _00377_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] VGND VGND VPWR
+ VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _04242_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or2_1
Xhold393 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] VGND VGND VPWR
+ VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
X_12951_ _05930_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _05931_ sky130_fd_sc_hd__nor2_1
X_11902_ _05028_ _05029_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__nand2_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _05862_
+ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ clknet_leaf_60_i_clk _00166_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11833_ _04966_ _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__nand2_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ clknet_leaf_35_i_clk _00098_ VGND VGND VPWR VPWR diff1\[11\] sky130_fd_sc_hd__dfxtp_1
X_11764_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] _04906_ VGND
+ VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__or4_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _03996_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__buf_2
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ clknet_leaf_25_i_clk _00029_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_1
X_11695_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04842_ VGND
+ VGND VPWR VPWR _04844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13434_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _06337_ VGND
+ VGND VPWR VPWR _06350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xrebuffer5 _04632_ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13365_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _06288_
+ _06216_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__a21o_1
X_10577_ _03872_ _03873_ _03874_ _03631_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15104_ clknet_leaf_115_i_clk _00649_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_1
X_12316_ _05383_ _05385_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13296_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _06230_
+ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__and2_1
X_15035_ clknet_leaf_92_i_clk _00580_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12247_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _05291_ VGND
+ VGND VPWR VPWR _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12178_ _05263_ _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__or2_4
X_11129_ _04012_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _04358_
+ _04359_ _04360_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14819_ clknet_leaf_75_i_clk _00364_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.valid_out
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_47_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08340_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[6\] _01900_ _01901_
+ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08271_ _01750_ _01840_ _01719_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07986_ net33 net51 VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__or2b_2
X_09725_ _02771_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09656_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _01876_ net273 _01945_ _02138_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _03006_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__mux2_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08538_ _02061_ _02073_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08469_ _02011_ _02012_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10500_ _03803_ _03804_ _03807_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11480_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _04662_ VGND
+ VGND VPWR VPWR _04663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10431_ net117 _03719_ _03744_ _03280_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13150_ _06093_ _06097_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__a21oi_1
X_10362_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[7\] _03681_ VGND
+ VGND VPWR VPWR _03682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12101_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _05191_
+ _05164_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13081_ _06037_ _06040_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__o21ai_1
X_10293_ _03623_ net252 _03620_ _03624_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__o211a_1
X_12032_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05139_ sky130_fd_sc_hd__buf_2
Xhold190 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND
+ VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13983_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06824_ _06553_
+ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__mux2_1
X_12934_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _05904_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12865_ _05857_ _05858_ _05567_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a21oi_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ clknet_leaf_45_i_clk _00149_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11816_ _04952_ _04930_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _05501_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] _05802_
+ _05803_ _05751_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ clknet_leaf_39_i_clk _00081_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11747_ _04850_ _04891_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14466_ clknet_leaf_39_i_clk _00012_ VGND VGND VPWR VPWR r_i_alpha1\[16\] sky130_fd_sc_hd__dfxtp_1
X_11678_ _04765_ _04829_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13417_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _05927_ VGND
+ VGND VPWR VPWR _06335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10629_ _03708_ _03922_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nor2_1
X_14397_ _07059_ _07177_ _07178_ _01475_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13348_ _06268_ _06270_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13279_ _05928_ _06213_ _06214_ _06216_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__a31o_1
X_15018_ clknet_leaf_95_i_clk _00563_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07840_ _01454_ net292 _01460_ _01462_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__o211a_1
X_07771_ net450 net3 _01411_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__mux2_1
X_09510_ _02844_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _02935_
+ _02936_ _02827_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__o221a_1
X_09441_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02873_ VGND
+ VGND VPWR VPWR _02874_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09372_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02814_
+ _02751_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08323_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\] VGND VGND VPWR VPWR _01887_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_145_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08254_ _01691_ _01830_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08185_ _01747_ _01762_ _01770_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07969_ _01565_ _01571_ _01572_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__a21oi_1
X_09708_ _03110_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__xnor2_1
X_10980_ _04011_ net419 _04219_ _04225_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__o211a_1
X_09639_ _03051_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12650_ _04455_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11601_ _04756_ net134 _04762_ _04766_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12581_ _05610_ _05611_ _05490_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14320_ _06909_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] VGND
+ VGND VPWR VPWR _07112_ sky130_fd_sc_hd__or2_1
X_11532_ _04707_ _04709_ _04376_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14251_ _07044_ _07047_ _07051_ _06926_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11463_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ net652 _04413_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__o31a_1
X_13202_ _06069_ _06153_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__and2_1
X_10414_ _03605_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _03728_
+ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__a22o_1
X_14182_ _06991_ _06992_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__or2b_1
X_11394_ _04579_ _04582_ _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a21oi_1
X_13133_ _06091_ _01512_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__and2b_1
X_10345_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _03664_
+ _03663_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _05998_ _06030_ _06031_ _05938_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__o211a_1
X_10276_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] _03609_
+ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__or2_1
X_12015_ _05128_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13966_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _06808_ VGND
+ VGND VPWR VPWR _06810_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12917_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05901_
+ _05842_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13897_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ _06716_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12848_ _03619_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__clkbuf_4
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12779_ _05781_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__clkbuf_4
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14518_ clknet_leaf_32_i_clk _00064_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14449_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _07157_ _07216_
+ _07219_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _03359_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08941_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[2\] _02341_ VGND VGND VPWR
+ VPWR _02431_ sky130_fd_sc_hd__o31a_1
X_08872_ _02371_ _02372_ _02344_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__mux2_1
X_07823_ _01333_ _01448_ _01449_ _01450_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07754_ _01402_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07685_ net20 _01350_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__or2_1
X_09424_ _02854_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09355_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _02796_
+ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08306_ net147 _01873_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__or2_1
X_09286_ _02329_ _02742_ _02743_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08237_ _01465_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08168_ _01757_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08099_ _01672_ _01654_ _01665_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__a21o_1
X_10130_ _03375_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10061_ _03425_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13820_ _06292_ _06680_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13751_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _06622_
+ _06562_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__o21ai_1
X_10963_ _04211_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12702_ _05715_ _05717_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__o21a_1
X_13682_ _06561_ net403 _06485_ _06564_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10894_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\]
+ _04132_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15421_ clknet_leaf_23_i_clk _00966_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12633_ _05485_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] VGND
+ VGND VPWR VPWR _05660_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15352_ clknet_leaf_29_i_clk _00897_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12564_ _05591_ _05593_ _05590_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a21o_1
X_14303_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _07042_ _07093_
+ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11515_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _04694_ VGND
+ VGND VPWR VPWR _04695_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15283_ clknet_leaf_16_i_clk _00828_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12495_ _05500_ net602 _05495_ _05538_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14234_ _06907_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _07038_ sky130_fd_sc_hd__or2_1
X_11446_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[8\] CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__or4_4
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14165_ _06646_ _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__nand2_1
X_11377_ _04444_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _04573_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13116_ _06070_ _06067_ _06074_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__or3b_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\] VGND VGND
+ VPWR VPWR _03654_ sky130_fd_sc_hd__inv_2
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _06915_ _06919_ _06904_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__a21o_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] _06003_ VGND
+ VGND VPWR VPWR _06017_ sky130_fd_sc_hd__xnor2_1
X_10259_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _03237_ _03601_
+ _03602_ _03258_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ clknet_leaf_109_i_clk _00543_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13949_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _06794_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07470_ _01095_ net452 _01194_ _01195_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09140_ _02607_ _02610_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09071_ _02313_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02548_
+ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08022_ _01472_ _01621_ _01464_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09973_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _03343_ VGND
+ VGND VPWR VPWR _03345_ sky130_fd_sc_hd__or2b_1
X_08924_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] _02415_ VGND
+ VGND VPWR VPWR _02416_ sky130_fd_sc_hd__xnor2_1
X_08855_ _02329_ net582 _02357_ _02358_ _02309_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__o221a_1
X_07806_ _01438_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08786_ _02300_ _02292_ _02294_ _02295_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__or4_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ net19 net20 _01385_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__and3_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07668_ _01338_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09407_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ _02836_ _02772_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07599_ diff2\[6\] _01270_ _01272_ diff3\[6\] _01284_ VGND VGND VPWR VPWR _01285_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09338_ _02785_ _02782_ _02784_ _02761_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09269_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _02726_ _02727_
+ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11300_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[13\] _04501_ VGND
+ VGND VPWR VPWR _04502_ sky130_fd_sc_hd__xnor2_1
X_12280_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[10\] CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ _05164_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11231_ _04379_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11162_ net134 _04379_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__or2_1
X_10113_ _03470_ _03460_ _03457_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__a21o_1
X_11093_ _04327_ _04328_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__and2_1
X_14921_ clknet_leaf_87_i_clk _00466_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_10044_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__buf_2
Xhold50 CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\] VGND VGND
+ VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 r_i_alpha1\[17\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 diff3\[4\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ clknet_4_6_0_i_clk _00397_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold83 diff3\[13\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _00309_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _06554_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _06665_
+ _06666_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__a22oi_1
X_14783_ clknet_leaf_74_i_clk _00328_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11995_ _05111_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__and2_1
X_13734_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _06606_
+ _06607_ _06584_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__o31ai_1
X_10946_ _04010_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] VGND
+ VGND VPWR VPWR _04197_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13665_ _06205_ _01979_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__and2_1
X_10877_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _04133_ VGND
+ VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12616_ _05643_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__nor2_1
X_15404_ clknet_leaf_34_i_clk _00949_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_13596_ _06491_ _06486_ _06487_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15335_ clknet_leaf_29_i_clk _00880_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12547_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _05573_ VGND
+ VGND VPWR VPWR _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15266_ clknet_leaf_10_i_clk _00811_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12478_ _05522_ _05523_ _05203_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14217_ _07021_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__clkbuf_4
X_11429_ _04613_ _04615_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__o21a_1
X_15197_ clknet_leaf_0_i_clk _00742_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14148_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06963_
+ _01862_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ _01861_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__clkbuf_4
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08640_ _02168_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08571_ _02103_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07522_ net69 net303 _01013_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__mux2_1
X_07453_ _01032_ _01085_ _01015_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_121_i_clk clknet_4_1_0_i_clk VGND VGND VPWR VPWR clknet_leaf_121_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07384_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ _01108_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09123_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[3\] VGND VGND VPWR
+ VPWR _02595_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09054_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _02525_ _02343_
+ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08005_ _01602_ _01605_ _01470_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold520 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] VGND VGND
+ VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\] VGND
+ VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09956_ _03191_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08907_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _02401_
+ _02320_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__o21ai_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _03264_ _03268_ _03183_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__a21o_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__clkbuf_4
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _02282_ _02285_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__xnor2_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _04064_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND
+ VGND VPWR VPWR _04065_ sky130_fd_sc_hd__nor2_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _04920_ _04921_ _04771_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__o21ai_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10731_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] _03999_
+ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13450_ _06356_ _06361_ _06364_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10662_ _03606_ _03952_ _03953_ _03780_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12401_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05423_ VGND
+ VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13381_ _06202_ _06301_ _06302_ _06110_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__o211a_1
X_10593_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03889_ VGND
+ VGND VPWR VPWR _03890_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15120_ clknet_leaf_116_i_clk _00665_ VGND VGND VPWR VPWR CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12332_ _05290_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15051_ clknet_leaf_111_i_clk net152 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12263_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[17\] _05291_ VGND
+ VGND VPWR VPWR _05340_ sky130_fd_sc_hd__xnor2_1
X_14002_ _06561_ net462 _06678_ _06841_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__o211a_1
X_11214_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _04420_
+ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__nand2_1
X_12194_ _05275_ _05276_ _05279_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput62 net62 VGND VGND VPWR VPWR out_alpha[13] sky130_fd_sc_hd__clkbuf_4
X_11145_ _04373_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
Xoutput73 net73 VGND VGND VPWR VPWR out_alpha[7] sky130_fd_sc_hd__clkbuf_4
Xoutput84 net84 VGND VGND VPWR VPWR out_costheta[17] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 VGND VGND VPWR VPWR out_sintheta[10] sky130_fd_sc_hd__clkbuf_4
X_11076_ _04205_ _04281_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__or2_1
X_14904_ clknet_leaf_87_i_clk _00449_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_10027_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] _03393_ VGND
+ VGND VPWR VPWR _03394_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14835_ clknet_leaf_77_i_clk _00380_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11978_ _05092_ _05095_ _05094_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14766_ clknet_leaf_51_i_clk _00311_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10929_ _04179_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__and2_1
X_13717_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _06580_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14697_ clknet_leaf_63_i_clk _00242_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13648_ _06535_ _06536_ _06205_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13579_ _06069_ _06477_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_i_clk clknet_4_12_0_i_clk VGND VGND VPWR VPWR clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15318_ clknet_leaf_22_i_clk _00863_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15249_ clknet_leaf_3_i_clk _00794_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_i_clk clknet_4_13_0_i_clk VGND VGND VPWR VPWR clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09810_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[2\] CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[1\]
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\] VGND VGND VPWR
+ VPWR _03204_ sky130_fd_sc_hd__and3_1
X_09741_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] _03144_ _03145_
+ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__a21o_1
X_09672_ _03081_ _03082_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__and2_2
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08623_ _01868_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[13\] VGND VGND VPWR VPWR
+ _02091_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07505_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _01159_ _01220_
+ _01221_ _01030_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__o221a_1
X_08485_ _02024_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07436_ _01044_ net193 _01169_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07367_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] _01099_ VGND
+ VGND VPWR VPWR _01108_ sky130_fd_sc_hd__or2_4
XFILLER_0_134_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09106_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _02579_ VGND
+ VGND VPWR VPWR _02580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07298_ _01026_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09037_ _02387_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _02517_
+ _02518_ _02414_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold350 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] VGND VGND
+ VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] VGND VGND
+ VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND VPWR VPWR
+ net500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold394 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[7\] VGND VGND VPWR VPWR
+ net511 sky130_fd_sc_hd__dlygate4sd3_1
X_09939_ _03306_ _03310_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__or2_1
X_12950_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_x\[11\] VGND VGND
+ VPWR VPWR _05930_ sky130_fd_sc_hd__inv_2
X_11901_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[5\] _05027_ VGND
+ VGND VPWR VPWR _05029_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12881_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ _05858_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__or3_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] _04930_ VGND
+ VGND VPWR VPWR _04967_ sky130_fd_sc_hd__nand2_1
X_14620_ clknet_leaf_58_i_clk _00165_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ clknet_leaf_35_i_clk _00097_ VGND VGND VPWR VPWR diff1\[10\] sky130_fd_sc_hd__dfxtp_1
X_11763_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _04905_ VGND
+ VGND VPWR VPWR _04906_ sky130_fd_sc_hd__xor2_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _03995_ net283 _03620_ _03998_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__o211a_1
X_13502_ _06216_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[16\] VGND
+ VGND VPWR VPWR _06409_ sky130_fd_sc_hd__and2_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ clknet_leaf_25_i_clk _00028_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11694_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[2\] _04842_ VGND
+ VGND VPWR VPWR _04843_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13433_ _06349_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10645_ _03923_ _03930_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13364_ net467 _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer6 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND VGND
+ VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_51_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10576_ _03872_ _03873_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a21oi_1
X_15103_ clknet_leaf_119_i_clk _00648_ VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12315_ _05383_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13295_ _06228_ _06229_ _05927_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15034_ clknet_leaf_97_i_clk _00579_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12246_ _05325_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__clkbuf_1
X_12177_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] _05262_ VGND
+ VGND VPWR VPWR _05264_ sky130_fd_sc_hd__nor2_1
X_11128_ _02308_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11059_ _04291_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14818_ clknet_leaf_74_i_clk _00363_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14749_ clknet_leaf_72_i_clk _00294_ VGND VGND VPWR VPWR CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08270_ _01843_ _01844_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07985_ net51 net33 VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__or2b_1
X_09724_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[13\]
+ _03107_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__or3_1
X_09655_ _03062_ _03064_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08606_ _02136_ _02137_ _01877_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _03001_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__xnor2_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _02022_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _02074_
+ _02075_ _02055_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08468_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[6\] _02010_ VGND VGND VPWR
+ VPWR _02012_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07419_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _01146_ VGND
+ VGND VPWR VPWR _01154_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08399_ _01876_ net427 _01945_ _01951_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10430_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ _03680_ _03671_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12100_ _05153_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ _05195_ _05196_ _05170_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13080_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06010_ VGND
+ VGND VPWR VPWR _06045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10292_ _03609_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\]
+ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12031_ _05130_ net201 _04979_ _05138_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__o211a_1
Xhold180 CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_x\[0\] VGND VGND VPWR
+ VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _00198_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
X_13982_ _06822_ _06823_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__xnor2_1
X_12933_ _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\]
+ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__or2_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ clknet_leaf_47_i_clk _00148_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11815_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[13\] CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[12\]
+ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__nor2_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _05800_ _05801_ _05490_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__o21ai_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _04754_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_y\[6\] _04889_
+ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__a22o_1
X_14534_ clknet_leaf_38_i_clk _00080_ VGND VGND VPWR VPWR CORDIC_PE\[0\].genblk1.cordic_engine_inst.in_alpha\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11677_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] VGND VGND
+ VPWR VPWR _04829_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14465_ clknet_leaf_38_i_clk _00011_ VGND VGND VPWR VPWR r_i_alpha1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13416_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__or2_1
X_10628_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _03921_ VGND
+ VGND VPWR VPWR _03922_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14396_ _06909_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND
+ VGND VPWR VPWR _07178_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13347_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06269_
+ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__nand2_1
X_10559_ _03848_ _03850_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13278_ _06200_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15017_ clknet_leaf_93_i_clk _00562_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12229_ _05307_ _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07770_ _01414_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
X_09440_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _02872_ VGND
+ VGND VPWR VPWR _02873_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09371_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _02814_
+ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08322_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[3\] CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[2\]
+ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND VPWR VPWR _01886_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08253_ _01700_ _01819_ _01829_ _01701_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_46_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08184_ _01747_ _01762_ _01770_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07968_ _01328_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__buf_4
X_09707_ _03100_ _03111_ _03114_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__o21a_1
X_07899_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_4
X_09638_ _03047_ _03050_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__and2_1
X_09569_ _02746_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _02989_
+ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11600_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[3\] _04765_
+ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12580_ _05610_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11531_ _04707_ _04709_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14250_ _07044_ _07047_ _07051_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11462_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] VGND VGND VPWR
+ VPWR _04646_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13201_ _05860_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[10\] _06151_
+ _06152_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__a22o_1
X_10413_ _03724_ _03727_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__o21a_1
X_14181_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[14\]
+ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] _06978_ _06934_
+ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__a41o_1
X_11393_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _04545_ VGND
+ VGND VPWR VPWR _04586_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13132_ _05844_ _06080_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__o21a_1
X_10344_ _03626_ net444 _03666_ _03667_ _03633_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _05853_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[12\] VGND
+ VGND VPWR VPWR _06031_ sky130_fd_sc_hd__or2_1
X_10275_ _03607_ net136 _03568_ _03613_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__o211a_1
X_12014_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.valid_out VGND VGND VPWR
+ VPWR _05128_ sky130_fd_sc_hd__inv_2
X_13965_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[4\] _06808_ VGND
+ VGND VPWR VPWR _06809_ sky130_fd_sc_hd__and2_1
X_12916_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] _05901_
+ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__nor2_1
X_13896_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[14\] _06707_ VGND
+ VGND VPWR VPWR _06748_ sky130_fd_sc_hd__xor2_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12847_ _05843_ net281 _05495_ _05846_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__o211a_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _05786_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14517_ clknet_leaf_33_i_clk _00063_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_1
X_11729_ _04874_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_y\[5\] VGND
+ VGND VPWR VPWR _04875_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14448_ _07222_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14379_ _06903_ CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _07162_
+ _07163_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08940_ _02430_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08871_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] _02365_
+ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__nand2_1
X_07822_ net361 _01344_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__and2_1
X_07753_ net418 _01401_ _01358_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__mux2_1
X_07684_ _01352_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09423_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] _02857_ VGND
+ VGND VPWR VPWR _02858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09354_ CORDIC_PE\[2\].genblk1.genblk1.cordic_engine_inst.out_alpha\[7\] _02794_
+ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08305_ _01868_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09285_ net626 _02320_ _01794_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08236_ _01656_ _01815_ _01329_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08167_ _01728_ _01756_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08098_ _01679_ _01680_ _01638_ _01672_ _01669_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_113_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10060_ _03024_ _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10962_ _03976_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__and2_1
X_13750_ _06292_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _06616_ _06621_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__o31a_1
X_12701_ _05715_ _05717_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10893_ _04023_ net118 _04147_ _04148_ _04059_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__o221a_1
X_13681_ _06563_ net453 VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ clknet_leaf_24_i_clk _00965_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_y\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12632_ _05657_ _05653_ _05654_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__or3_1
XFILLER_0_81_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12563_ _05596_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
X_15351_ clknet_leaf_47_i_clk _00896_ VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11514_ _04692_ _04693_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__or2b_4
X_14302_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[15\] _07041_ VGND
+ VGND VPWR VPWR _07096_ sky130_fd_sc_hd__xnor2_1
X_12494_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\] _05536_
+ _05537_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__a21o_1
X_15282_ clknet_leaf_51_i_clk _00827_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11445_ _04623_ _04625_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__a21oi_2
X_14233_ _07035_ _07036_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14164_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\] CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ _06967_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11376_ _04570_ _04571_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ _06070_ _06067_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__o21bai_2
X_10327_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ _03634_ _03651_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14095_ _06915_ _06919_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__nor2_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[9\] _06010_ _06005_
+ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__o21ai_1
X_10258_ _03599_ _03600_ _03201_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10189_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[8\] _03523_ _03530_
+ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[9\] VGND VGND VPWR VPWR
+ _03540_ sky130_fd_sc_hd__a22o_1
X_14997_ clknet_leaf_108_i_clk _00542_ VGND VGND VPWR VPWR CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13948_ _06793_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13879_ _06556_ _06731_ _06733_ _06459_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09070_ _02542_ _02547_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08021_ _01612_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09972_ _03343_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_y\[7\] VGND
+ VGND VPWR VPWR _03344_ sky130_fd_sc_hd__or2b_1
X_08923_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\] CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[2\]
+ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08854_ _02356_ _02354_ _02355_ _02320_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__o31ai_1
X_07805_ net382 _01437_ _01411_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08785_ _02292_ _02294_ _02295_ _02300_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__o31a_1
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ net199 _01345_ _01388_ _01389_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__a22o_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07667_ _00991_ _01334_ net16 VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09406_ _02750_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07598_ _01273_ diff1\[6\] VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09337_ _02782_ _02784_ _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09268_ _02726_ _02727_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[15\]
+ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08219_ _01598_ _01612_ _01800_ _01470_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_09199_ _02657_ _02649_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__and2b_1
X_11230_ CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_alpha\[16\] _04439_
+ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__xnor2_1
X_11161_ _04377_ net222 _04219_ _04384_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10112_ _03031_ _03455_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__nand2_1
X_11092_ _04325_ _04326_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[11\]
+ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__o21ai_2
X_14920_ clknet_leaf_83_i_clk _00465_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10043_ _03407_ _03408_ _03207_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__mux2_1
Xhold40 CORDIC_PE\[6\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND VGND
+ VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 net106 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\] VGND VGND
+ VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ clknet_4_7_0_i_clk _00396_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold73 diff1\[7\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] VGND VGND
+ VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[0\] VGND
+ VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _06658_ _06659_ _06664_ _06553_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__o31a_1
X_14782_ clknet_leaf_76_i_clk _00327_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_11994_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_x\[15\] _05081_ VGND
+ VGND VPWR VPWR _05112_ sky130_fd_sc_hd__xor2_1
X_13733_ _06606_ _06607_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\]
+ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__o21a_1
X_10945_ _04194_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13664_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[17\] _06210_ _06550_
+ _06551_ _06526_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10876_ _04108_ _04132_ _04035_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__o21ai_1
X_15403_ clknet_leaf_31_i_clk _00948_ VGND VGND VPWR VPWR CORDIC_PE\[14\].genblk1.genblk1.cordic_engine_inst.out_alpha\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12615_ _05642_ _05636_ _05638_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13595_ _06486_ _06487_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__a21oi_1
X_15334_ clknet_leaf_23_i_clk net221 VGND VGND VPWR VPWR CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_quadrant\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12546_ _05579_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15265_ clknet_leaf_10_i_clk _00810_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_x\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[8\] _05516_
+ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_alpha\[9\] VGND VGND VPWR
+ VPWR _05523_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14216_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_y\[3\] _07019_ _07021_
+ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11428_ _04613_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__nand2_1
X_15196_ clknet_leaf_0_i_clk _00741_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_y\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11359_ _04556_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14147_ CORDIC_PE\[13\].genblk1.genblk1.cordic_engine_inst.out_alpha\[10\] _06963_
+ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ _06905_ net256 _06678_ _06906_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__o211a_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _05966_ _05973_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2_1
X_08570_ _02082_ _02088_ _02095_ _02105_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__o31ai_2
X_07521_ _01232_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07452_ _01076_ _01040_ _01181_ _01085_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_07383_ _01037_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09122_ _02594_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09053_ _02530_ _02524_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_08004_ _01603_ _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold510 CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\] VGND VGND
+ VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold521 CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[4\] VGND VGND VPWR VPWR
+ net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_y\[0\] VGND VGND VPWR
+ VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09955_ _03327_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__xnor2_1
X_08906_ CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\] _02401_
+ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__and2_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _03264_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nor2_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__buf_2
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_y\[16\] _02284_ VGND VGND VPWR
+ VPWR _02285_ sky130_fd_sc_hd__xor2_2
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _01377_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08699_ CORDIC_PE\[0\].genblk1.cordic_engine_inst.out_x\[9\] _02221_ VGND VGND VPWR
+ VPWR _02222_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10730_ _03995_ net179 _04003_ _04007_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_10661_ _03608_ CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_x\[12\] VGND
+ VGND VPWR VPWR _03953_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12400_ CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_x\[14\] _05423_ VGND
+ VGND VPWR VPWR _05462_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13380_ _06251_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_y\[1\] VGND
+ VGND VPWR VPWR _06302_ sky130_fd_sc_hd__or2_1
X_10592_ CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_y\[11\] _03650_ _03880_
+ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_12331_ CORDIC_PE\[9\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _05400_ _01249_
+ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12262_ _05332_ _05335_ _05331_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__o21ai_1
X_15050_ clknet_leaf_110_i_clk net123 VGND VGND VPWR VPWR CORDIC_PE\[8\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_11213_ _04390_ CORDIC_PE\[7\].genblk1.genblk1.cordic_engine_inst.out_alpha\[13\]
+ _04387_ _04425_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__o211a_1
X_14001_ _06839_ _06840_ _06584_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__o21ai_1
X_12193_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__clkbuf_4
X_11144_ _03997_ _02310_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and2_1
Xoutput63 net63 VGND VGND VPWR VPWR out_alpha[14] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR out_alpha[8] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 VGND VGND VPWR VPWR out_costheta[1] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 VGND VGND VPWR VPWR out_sintheta[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11075_ _04310_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__nand2_1
X_14903_ clknet_leaf_87_i_clk _00448_ VGND VGND VPWR VPWR CORDIC_PE\[5\].genblk1.genblk1.cordic_engine_inst.out_y\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_10026_ CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_x\[16\] _03392_ VGND
+ VGND VPWR VPWR _03393_ sky130_fd_sc_hd__xnor2_1
X_14834_ clknet_leaf_77_i_clk _00379_ VGND VGND VPWR VPWR CORDIC_PE\[4\].genblk1.genblk1.cordic_engine_inst.out_alpha\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14765_ clknet_leaf_16_i_clk _00310_ VGND VGND VPWR VPWR CORDIC_PE\[3\].genblk1.genblk1.cordic_engine_inst.out_alpha\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11977_ _04862_ _05096_ _05097_ _05080_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13716_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[6\] CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[5\]
+ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_alpha\[4\] _06571_ VGND VGND
+ VPWR VPWR _06593_ sky130_fd_sc_hd__and4_1
X_10928_ _04178_ _04180_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_14696_ clknet_leaf_61_i_clk _00241_ VGND VGND VPWR VPWR CORDIC_PE\[1\].genblk1.genblk1.cordic_engine_inst.out_x\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_13647_ _06535_ _06536_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__and2_1
X_10859_ _03976_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[6\] _06476_ CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.valid_out
+ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_15317_ clknet_leaf_23_i_clk _00862_ VGND VGND VPWR VPWR CORDIC_PE\[12\].genblk1.genblk1.cordic_engine_inst.out_x\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12529_ _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__buf_2
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15248_ clknet_leaf_8_i_clk _00793_ VGND VGND VPWR VPWR CORDIC_PE\[11\].genblk1.genblk1.cordic_engine_inst.out_y\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15179_ clknet_leaf_115_i_clk _00724_ VGND VGND VPWR VPWR CORDIC_PE\[10\].genblk1.genblk1.cordic_engine_inst.out_alpha\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09740_ _03133_ _03138_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__and2b_1
.ends

