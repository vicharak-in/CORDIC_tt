VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cordic_tt_top
  CLASS BLOCK ;
  FOREIGN cordic_tt_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 442.310 BY 453.030 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 10.640 16.620 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.620 10.640 170.220 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 322.220 10.640 323.820 440.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.380 436.780 21.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 173.560 436.780 175.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.740 436.780 328.340 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.320 10.640 166.920 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 318.920 10.640 320.520 440.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.080 436.780 18.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 170.260 436.780 171.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 323.440 436.780 325.040 ;
    END
  END VPWR
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 438.310 225.800 442.310 226.400 ;
    END
  END i_clk
  PIN i_rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END i_rst_n
  PIN i_valid_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END i_valid_in
  PIN in_alpha[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 154.190 449.030 154.470 453.030 ;
    END
  END in_alpha[0]
  PIN in_alpha[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 232.390 449.030 232.670 453.030 ;
    END
  END in_alpha[10]
  PIN in_alpha[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 449.030 240.490 453.030 ;
    END
  END in_alpha[11]
  PIN in_alpha[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 449.030 248.310 453.030 ;
    END
  END in_alpha[12]
  PIN in_alpha[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 255.850 449.030 256.130 453.030 ;
    END
  END in_alpha[13]
  PIN in_alpha[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 263.670 449.030 263.950 453.030 ;
    END
  END in_alpha[14]
  PIN in_alpha[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 271.490 449.030 271.770 453.030 ;
    END
  END in_alpha[15]
  PIN in_alpha[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 279.310 449.030 279.590 453.030 ;
    END
  END in_alpha[16]
  PIN in_alpha[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 287.130 449.030 287.410 453.030 ;
    END
  END in_alpha[17]
  PIN in_alpha[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 162.010 449.030 162.290 453.030 ;
    END
  END in_alpha[1]
  PIN in_alpha[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 169.830 449.030 170.110 453.030 ;
    END
  END in_alpha[2]
  PIN in_alpha[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.650 449.030 177.930 453.030 ;
    END
  END in_alpha[3]
  PIN in_alpha[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.470 449.030 185.750 453.030 ;
    END
  END in_alpha[4]
  PIN in_alpha[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 449.030 193.570 453.030 ;
    END
  END in_alpha[5]
  PIN in_alpha[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 201.110 449.030 201.390 453.030 ;
    END
  END in_alpha[6]
  PIN in_alpha[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 208.930 449.030 209.210 453.030 ;
    END
  END in_alpha[7]
  PIN in_alpha[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 216.750 449.030 217.030 453.030 ;
    END
  END in_alpha[8]
  PIN in_alpha[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 224.570 449.030 224.850 453.030 ;
    END
  END in_alpha[9]
  PIN in_x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 13.430 449.030 13.710 453.030 ;
    END
  END in_x[0]
  PIN in_x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 91.630 449.030 91.910 453.030 ;
    END
  END in_x[10]
  PIN in_x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 449.030 99.730 453.030 ;
    END
  END in_x[11]
  PIN in_x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 449.030 107.550 453.030 ;
    END
  END in_x[12]
  PIN in_x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 449.030 115.370 453.030 ;
    END
  END in_x[13]
  PIN in_x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 122.910 449.030 123.190 453.030 ;
    END
  END in_x[14]
  PIN in_x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 130.730 449.030 131.010 453.030 ;
    END
  END in_x[15]
  PIN in_x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 449.030 138.830 453.030 ;
    END
  END in_x[16]
  PIN in_x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.370 449.030 146.650 453.030 ;
    END
  END in_x[17]
  PIN in_x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 21.250 449.030 21.530 453.030 ;
    END
  END in_x[1]
  PIN in_x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 449.030 29.350 453.030 ;
    END
  END in_x[2]
  PIN in_x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 449.030 37.170 453.030 ;
    END
  END in_x[3]
  PIN in_x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 44.710 449.030 44.990 453.030 ;
    END
  END in_x[4]
  PIN in_x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.530 449.030 52.810 453.030 ;
    END
  END in_x[5]
  PIN in_x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 60.350 449.030 60.630 453.030 ;
    END
  END in_x[6]
  PIN in_x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 449.030 68.450 453.030 ;
    END
  END in_x[7]
  PIN in_x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 75.990 449.030 76.270 453.030 ;
    END
  END in_x[8]
  PIN in_x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 449.030 84.090 453.030 ;
    END
  END in_x[9]
  PIN in_y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 294.950 449.030 295.230 453.030 ;
    END
  END in_y[0]
  PIN in_y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 373.150 449.030 373.430 453.030 ;
    END
  END in_y[10]
  PIN in_y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 380.970 449.030 381.250 453.030 ;
    END
  END in_y[11]
  PIN in_y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 388.790 449.030 389.070 453.030 ;
    END
  END in_y[12]
  PIN in_y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 396.610 449.030 396.890 453.030 ;
    END
  END in_y[13]
  PIN in_y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 404.430 449.030 404.710 453.030 ;
    END
  END in_y[14]
  PIN in_y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 449.030 412.530 453.030 ;
    END
  END in_y[15]
  PIN in_y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 420.070 449.030 420.350 453.030 ;
    END
  END in_y[16]
  PIN in_y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 427.890 449.030 428.170 453.030 ;
    END
  END in_y[17]
  PIN in_y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 449.030 303.050 453.030 ;
    END
  END in_y[1]
  PIN in_y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 310.590 449.030 310.870 453.030 ;
    END
  END in_y[2]
  PIN in_y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 449.030 318.690 453.030 ;
    END
  END in_y[3]
  PIN in_y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 326.230 449.030 326.510 453.030 ;
    END
  END in_y[4]
  PIN in_y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 334.050 449.030 334.330 453.030 ;
    END
  END in_y[5]
  PIN in_y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 341.870 449.030 342.150 453.030 ;
    END
  END in_y[6]
  PIN in_y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 349.690 449.030 349.970 453.030 ;
    END
  END in_y[7]
  PIN in_y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 449.030 357.790 453.030 ;
    END
  END in_y[8]
  PIN in_y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 449.030 365.610 453.030 ;
    END
  END in_y[9]
  PIN o_valid_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END o_valid_out
  PIN out_alpha[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END out_alpha[0]
  PIN out_alpha[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END out_alpha[10]
  PIN out_alpha[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END out_alpha[11]
  PIN out_alpha[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END out_alpha[12]
  PIN out_alpha[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END out_alpha[13]
  PIN out_alpha[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END out_alpha[14]
  PIN out_alpha[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END out_alpha[15]
  PIN out_alpha[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END out_alpha[16]
  PIN out_alpha[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END out_alpha[17]
  PIN out_alpha[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END out_alpha[1]
  PIN out_alpha[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END out_alpha[2]
  PIN out_alpha[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END out_alpha[3]
  PIN out_alpha[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END out_alpha[4]
  PIN out_alpha[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END out_alpha[5]
  PIN out_alpha[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END out_alpha[6]
  PIN out_alpha[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END out_alpha[7]
  PIN out_alpha[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END out_alpha[8]
  PIN out_alpha[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END out_alpha[9]
  PIN out_costheta[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END out_costheta[0]
  PIN out_costheta[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END out_costheta[10]
  PIN out_costheta[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END out_costheta[11]
  PIN out_costheta[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END out_costheta[12]
  PIN out_costheta[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END out_costheta[13]
  PIN out_costheta[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END out_costheta[14]
  PIN out_costheta[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END out_costheta[15]
  PIN out_costheta[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END out_costheta[16]
  PIN out_costheta[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END out_costheta[17]
  PIN out_costheta[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END out_costheta[1]
  PIN out_costheta[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END out_costheta[2]
  PIN out_costheta[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END out_costheta[3]
  PIN out_costheta[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END out_costheta[4]
  PIN out_costheta[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END out_costheta[5]
  PIN out_costheta[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END out_costheta[6]
  PIN out_costheta[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END out_costheta[7]
  PIN out_costheta[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END out_costheta[8]
  PIN out_costheta[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END out_costheta[9]
  PIN out_sintheta[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END out_sintheta[0]
  PIN out_sintheta[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END out_sintheta[10]
  PIN out_sintheta[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END out_sintheta[11]
  PIN out_sintheta[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END out_sintheta[12]
  PIN out_sintheta[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END out_sintheta[13]
  PIN out_sintheta[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END out_sintheta[14]
  PIN out_sintheta[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END out_sintheta[15]
  PIN out_sintheta[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END out_sintheta[16]
  PIN out_sintheta[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END out_sintheta[17]
  PIN out_sintheta[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END out_sintheta[1]
  PIN out_sintheta[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END out_sintheta[2]
  PIN out_sintheta[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END out_sintheta[3]
  PIN out_sintheta[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END out_sintheta[4]
  PIN out_sintheta[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END out_sintheta[5]
  PIN out_sintheta[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END out_sintheta[6]
  PIN out_sintheta[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END out_sintheta[7]
  PIN out_sintheta[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END out_sintheta[8]
  PIN out_sintheta[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END out_sintheta[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 436.540 440.725 ;
      LAYER met1 ;
        RECT 4.670 10.640 436.540 444.680 ;
      LAYER met2 ;
        RECT 4.690 448.750 13.150 449.030 ;
        RECT 13.990 448.750 20.970 449.030 ;
        RECT 21.810 448.750 28.790 449.030 ;
        RECT 29.630 448.750 36.610 449.030 ;
        RECT 37.450 448.750 44.430 449.030 ;
        RECT 45.270 448.750 52.250 449.030 ;
        RECT 53.090 448.750 60.070 449.030 ;
        RECT 60.910 448.750 67.890 449.030 ;
        RECT 68.730 448.750 75.710 449.030 ;
        RECT 76.550 448.750 83.530 449.030 ;
        RECT 84.370 448.750 91.350 449.030 ;
        RECT 92.190 448.750 99.170 449.030 ;
        RECT 100.010 448.750 106.990 449.030 ;
        RECT 107.830 448.750 114.810 449.030 ;
        RECT 115.650 448.750 122.630 449.030 ;
        RECT 123.470 448.750 130.450 449.030 ;
        RECT 131.290 448.750 138.270 449.030 ;
        RECT 139.110 448.750 146.090 449.030 ;
        RECT 146.930 448.750 153.910 449.030 ;
        RECT 154.750 448.750 161.730 449.030 ;
        RECT 162.570 448.750 169.550 449.030 ;
        RECT 170.390 448.750 177.370 449.030 ;
        RECT 178.210 448.750 185.190 449.030 ;
        RECT 186.030 448.750 193.010 449.030 ;
        RECT 193.850 448.750 200.830 449.030 ;
        RECT 201.670 448.750 208.650 449.030 ;
        RECT 209.490 448.750 216.470 449.030 ;
        RECT 217.310 448.750 224.290 449.030 ;
        RECT 225.130 448.750 232.110 449.030 ;
        RECT 232.950 448.750 239.930 449.030 ;
        RECT 240.770 448.750 247.750 449.030 ;
        RECT 248.590 448.750 255.570 449.030 ;
        RECT 256.410 448.750 263.390 449.030 ;
        RECT 264.230 448.750 271.210 449.030 ;
        RECT 272.050 448.750 279.030 449.030 ;
        RECT 279.870 448.750 286.850 449.030 ;
        RECT 287.690 448.750 294.670 449.030 ;
        RECT 295.510 448.750 302.490 449.030 ;
        RECT 303.330 448.750 310.310 449.030 ;
        RECT 311.150 448.750 318.130 449.030 ;
        RECT 318.970 448.750 325.950 449.030 ;
        RECT 326.790 448.750 333.770 449.030 ;
        RECT 334.610 448.750 341.590 449.030 ;
        RECT 342.430 448.750 349.410 449.030 ;
        RECT 350.250 448.750 357.230 449.030 ;
        RECT 358.070 448.750 365.050 449.030 ;
        RECT 365.890 448.750 372.870 449.030 ;
        RECT 373.710 448.750 380.690 449.030 ;
        RECT 381.530 448.750 388.510 449.030 ;
        RECT 389.350 448.750 396.330 449.030 ;
        RECT 397.170 448.750 404.150 449.030 ;
        RECT 404.990 448.750 411.970 449.030 ;
        RECT 412.810 448.750 419.790 449.030 ;
        RECT 420.630 448.750 427.610 449.030 ;
        RECT 428.450 448.750 429.550 449.030 ;
        RECT 4.690 4.280 429.550 448.750 ;
        RECT 4.690 4.000 220.610 4.280 ;
        RECT 221.450 4.000 367.810 4.280 ;
        RECT 368.650 4.000 429.550 4.280 ;
      LAYER met3 ;
        RECT 4.400 445.720 438.310 446.570 ;
        RECT 3.990 438.960 438.310 445.720 ;
        RECT 4.400 437.560 438.310 438.960 ;
        RECT 3.990 430.800 438.310 437.560 ;
        RECT 4.400 429.400 438.310 430.800 ;
        RECT 3.990 422.640 438.310 429.400 ;
        RECT 4.400 421.240 438.310 422.640 ;
        RECT 3.990 414.480 438.310 421.240 ;
        RECT 4.400 413.080 438.310 414.480 ;
        RECT 3.990 406.320 438.310 413.080 ;
        RECT 4.400 404.920 438.310 406.320 ;
        RECT 3.990 398.160 438.310 404.920 ;
        RECT 4.400 396.760 438.310 398.160 ;
        RECT 3.990 390.000 438.310 396.760 ;
        RECT 4.400 388.600 438.310 390.000 ;
        RECT 3.990 381.840 438.310 388.600 ;
        RECT 4.400 380.440 438.310 381.840 ;
        RECT 3.990 373.680 438.310 380.440 ;
        RECT 4.400 372.280 438.310 373.680 ;
        RECT 3.990 365.520 438.310 372.280 ;
        RECT 4.400 364.120 438.310 365.520 ;
        RECT 3.990 357.360 438.310 364.120 ;
        RECT 4.400 355.960 438.310 357.360 ;
        RECT 3.990 349.200 438.310 355.960 ;
        RECT 4.400 347.800 438.310 349.200 ;
        RECT 3.990 341.040 438.310 347.800 ;
        RECT 4.400 339.640 438.310 341.040 ;
        RECT 3.990 332.880 438.310 339.640 ;
        RECT 4.400 331.480 438.310 332.880 ;
        RECT 3.990 324.720 438.310 331.480 ;
        RECT 4.400 323.320 438.310 324.720 ;
        RECT 3.990 316.560 438.310 323.320 ;
        RECT 4.400 315.160 438.310 316.560 ;
        RECT 3.990 308.400 438.310 315.160 ;
        RECT 4.400 307.000 438.310 308.400 ;
        RECT 3.990 300.240 438.310 307.000 ;
        RECT 4.400 298.840 438.310 300.240 ;
        RECT 3.990 292.080 438.310 298.840 ;
        RECT 4.400 290.680 438.310 292.080 ;
        RECT 3.990 283.920 438.310 290.680 ;
        RECT 4.400 282.520 438.310 283.920 ;
        RECT 3.990 275.760 438.310 282.520 ;
        RECT 4.400 274.360 438.310 275.760 ;
        RECT 3.990 267.600 438.310 274.360 ;
        RECT 4.400 266.200 438.310 267.600 ;
        RECT 3.990 259.440 438.310 266.200 ;
        RECT 4.400 258.040 438.310 259.440 ;
        RECT 3.990 251.280 438.310 258.040 ;
        RECT 4.400 249.880 438.310 251.280 ;
        RECT 3.990 243.120 438.310 249.880 ;
        RECT 4.400 241.720 438.310 243.120 ;
        RECT 3.990 234.960 438.310 241.720 ;
        RECT 4.400 233.560 438.310 234.960 ;
        RECT 3.990 226.800 438.310 233.560 ;
        RECT 4.400 225.400 437.910 226.800 ;
        RECT 3.990 218.640 438.310 225.400 ;
        RECT 4.400 217.240 438.310 218.640 ;
        RECT 3.990 210.480 438.310 217.240 ;
        RECT 4.400 209.080 438.310 210.480 ;
        RECT 3.990 202.320 438.310 209.080 ;
        RECT 4.400 200.920 438.310 202.320 ;
        RECT 3.990 194.160 438.310 200.920 ;
        RECT 4.400 192.760 438.310 194.160 ;
        RECT 3.990 186.000 438.310 192.760 ;
        RECT 4.400 184.600 438.310 186.000 ;
        RECT 3.990 177.840 438.310 184.600 ;
        RECT 4.400 176.440 438.310 177.840 ;
        RECT 3.990 169.680 438.310 176.440 ;
        RECT 4.400 168.280 438.310 169.680 ;
        RECT 3.990 161.520 438.310 168.280 ;
        RECT 4.400 160.120 438.310 161.520 ;
        RECT 3.990 153.360 438.310 160.120 ;
        RECT 4.400 151.960 438.310 153.360 ;
        RECT 3.990 145.200 438.310 151.960 ;
        RECT 4.400 143.800 438.310 145.200 ;
        RECT 3.990 137.040 438.310 143.800 ;
        RECT 4.400 135.640 438.310 137.040 ;
        RECT 3.990 128.880 438.310 135.640 ;
        RECT 4.400 127.480 438.310 128.880 ;
        RECT 3.990 120.720 438.310 127.480 ;
        RECT 4.400 119.320 438.310 120.720 ;
        RECT 3.990 112.560 438.310 119.320 ;
        RECT 4.400 111.160 438.310 112.560 ;
        RECT 3.990 104.400 438.310 111.160 ;
        RECT 4.400 103.000 438.310 104.400 ;
        RECT 3.990 96.240 438.310 103.000 ;
        RECT 4.400 94.840 438.310 96.240 ;
        RECT 3.990 88.080 438.310 94.840 ;
        RECT 4.400 86.680 438.310 88.080 ;
        RECT 3.990 79.920 438.310 86.680 ;
        RECT 4.400 78.520 438.310 79.920 ;
        RECT 3.990 71.760 438.310 78.520 ;
        RECT 4.400 70.360 438.310 71.760 ;
        RECT 3.990 63.600 438.310 70.360 ;
        RECT 4.400 62.200 438.310 63.600 ;
        RECT 3.990 55.440 438.310 62.200 ;
        RECT 4.400 54.040 438.310 55.440 ;
        RECT 3.990 47.280 438.310 54.040 ;
        RECT 4.400 45.880 438.310 47.280 ;
        RECT 3.990 39.120 438.310 45.880 ;
        RECT 4.400 37.720 438.310 39.120 ;
        RECT 3.990 30.960 438.310 37.720 ;
        RECT 4.400 29.560 438.310 30.960 ;
        RECT 3.990 22.800 438.310 29.560 ;
        RECT 4.400 21.400 438.310 22.800 ;
        RECT 3.990 14.640 438.310 21.400 ;
        RECT 4.400 13.240 438.310 14.640 ;
        RECT 3.990 6.480 438.310 13.240 ;
        RECT 4.400 5.630 438.310 6.480 ;
      LAYER met4 ;
        RECT 14.095 34.855 14.620 407.825 ;
        RECT 17.020 34.855 164.920 407.825 ;
        RECT 167.320 34.855 168.220 407.825 ;
        RECT 170.620 34.855 318.520 407.825 ;
        RECT 320.920 34.855 321.820 407.825 ;
        RECT 324.220 34.855 351.145 407.825 ;
  END
END cordic_tt_top
END LIBRARY

